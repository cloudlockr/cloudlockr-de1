��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�~Zڟe���!Db��>Y|s�_�=AX����N!��z��u����8�A��ԛ�VN�{CBr�������1}f���S9T�����M��8�e�RzSpW��ά��ɻ�+�Q�+R=�a^�HsR�9O��Tx���;'A�Wf/P��
��ȥmZB3R�/d�w����������L�@q�z�f����EX���9�(X�Fݝv�H�r�����TL'a��T�x-.cSE�qG�c��'��	n���2��\�F՜^	'��%\i�z��͸\r�2�2�Iq.��'�FP�� ���->Q	��o#2�~��AuHjC����|��"4 ��q�+���D�(X�������1\Šr�Af�:,f�f�;�dK�C)[J2��L4k~*2��Ђw-~a�zM��UO9�,�Ko+�8Շ�������xչX��wE���(�(�k�zu����i���i�D7L���!�g�o��P��4�j�$վ�: r/x=	��s�	U48'X�^�W�t�'�;XN����Gz����=do����~�X{��V���<j��^�mi��/=�`;H��@W�)2��2!�g./e��v��/g8-���+���Qm_�����%��!���������H�'���z5�P����;�/���٨�ju�<f_x�5�n4���_ �C�e=N�R�j��Ϧ ;�.ĭa_�O.�]0�o	��}D��𻑖�3 �B�]��	+�O�"�׊j�TP�e���汪�3'����'{i�f����$.�P\#�'zG��SUz�qjz��m\9"�ңS�����X;9����X���W�h�+
Iw��¶�.<�Y���?�Z�6�"�)аm��t3��D�̎,m�}�!��a�gxr��I4]��q��9�GG��Vϓ�P�?������UL%�<���n�������8��zʙS�(�A�H*N3	~������@��Iq`>ǃ-ܿ0���u)���f1�،��do�T��Hmk�ƹJ�Ӌ��y���7b���@�(�g��@�`a-���9j�E�2'B�y��;+8�n��@�	G��A��C'A'�Ev�F�qYE�C�R��)`Z�|e��1 +È�Z�\a�5��*��(SnE9���Lv0Fehv���u}��?��Zr��]0c�b 2j�Ł�
a��s��;�	��>p<�EN�J��Sf�Z�cT��8�>��
�D4�'� p�_Q#uXMʬ_:&����%�h�C7��2�X&���h�Ԭ���t�����ܺB/Idp���V�g�TO�m�����Dxɺ���n�&��s� p����~ٯ�?6�W�5E�O6�U�0=��,8Rjf��v��!R/�`5��ú�7Xf>spJNr|����o�(��ޒD�u�N!iQy�8<�ث"QE�=ð9�l��ŇV�dJA�fe��	�
'���sx��e�}�'I���1R�6���O�, �hL4YJ��~ɠ�N���0ٰ�8n�2lTL������Ǫ�AH�m�^�/X"�+��� �e�x�p�:��i���хP2���+�g6��f��딕TwS���]~�)YPeTq�P��U�u䬄]ȗ�	���^���
���ֵ�RM����R��o;-Ԃj�:Rw�/{{�9�3�*�T%Spy(��XK̀�S.9��CT�6�s�i��K���������7��s�#����a�^�{H�y�97���&��Lu�T�2�\�Jr��#��A�f�t����(0�w��u�T+A����`#�Dt�<&y9,ַ��L*�Z{��2E���A*��_���y#���6s�N�Q��L]��ޙFf2����9f��t�B�c�T�R}�a]��k
����%�K�eX�fiF��KFG�n�yՓwi̧�;vԠT�1���Ā|s�����_�0��N���X���tS��ժ@Zq=|�����li�Ye��k$�������/�$������1ߠs{�4`���.�FX�>xs��#��¬�梭-�j�ԓ��r��<(�U�U��Yu�yn��H��� ڷ�y���τ������E�W]���O؉c�x�?�)�+�=�׬D��%̅8Z��|�!�,��z��ycu�P�7��Ē>]+�]=�Kb�JXFh��@���,Ԟ�5��r��}�%r�C���#|�`c�����
`��c�P�eC�����.�Ci�|*�sIiErU���m8��wR	:��[�~��'�����s���SM��qA��zc���p_���޶ ѵ6�3r%P-�;`�{S�7J�D��T��p�m��#J��)����I�Σ6���<�"<t��6&$��Z�{Ư��Z��e�D�	"�pzF崪6vhsG�_�����<��b�6��]3x~7��*����k�����\gw���|�059h���h'te�� i  �ш�Ru��{����R+��=M>�N/��|P̥Q�I�pWZNa��ª�Zd�AQ� j�*��f�tY�{����"s�y2�����(��P��5��Y�RN�F����iy8��A�6�e�g�Ǻ3�!�30���r'�>n���;]e�e���e �R-uA�5�E�������4q����=AB}y�� D���� �  �oɆ��u2�J�YN"�z���ً( �P(�L�?���%��[<���K4A���p�a'2N����w�N�X���A����R9p��$�(��Ԫ}��2,zgV��lL��h6��.�v���Kp%��,���f�g�_}�J��T7S�h;?���Fn����ƌ�/wc/��0J��J��8�z��lK@�	�+W$�CW��ts���r�q�+�rnc=�]K)��f������1=��j�H�Ѡ|�r/en���Y[�E��c����N�q��Ӣ˺�[o�93Q2�Z���x��7���9�Qg�a`��R����h��=�@��7�(p�ؗRk8�M�3mé��H)�����*C�~;���`�q��.��̺n�K
�A�2r�R���S@?P��\(U�(���Rƴ=�6�#����5�cy-8�5��fL# �u�mi�> %l���/b�c�3��u���,L��?(�[1�N�sg2]� ��09Ojvz�8�4)�\e^��}�6�X+A��-@�?N�R���Rn[ ǔ���_�~�4bu�%�=H��,�3��d���Wxql>�ծ[����a|ȿ���h��2bi�'