��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�~Zڟe�ͤ3��5?��^~��Ha�ptƼⷞ\T���ҚO��'���v��rR���ϗ��Qv_A�Z*�	m3�̻:�J�ʟ'�*�)�A C�S�u�9cd�!YnQ�?��k��U�������J0�!3iˀDX��LYܪȉF)�ݜ"/�'�fÐ1�E��> s���^a�N.�Hc��c�ە��[�]!������ ��$�I�#�4.�R1�:���afu�7l�m5�{)���be;�aN���[ ��\�-+��%�r���)���\dV�D��#��{H�O��e�Vv��m�:n��q���졿�O'�Yz��!�*���> �?�	�մq�,������� B�^����bt9�o�t����hT,�h�&H&������~���f��*�e�L.:�(�_��s��ԛ��}��.�}��i'� -�\��4Su��C ���xn&�ˮ��<��������)�u�X����&v!N1|[0�c�R0j�0��Z8!=�|I�'|�t��]�h���A�.��t��k��Nj5${VA�UG�Iؿyb�q�g~�O�f�@+���*�`�Z�n~p^�����EJkl�������R��;[l\<\������:�}�z�!_?�4����G��U�o�_W���&�H��	�(X��0��iOM01��C�~e�i��V��ؓan��
�`A�:��j�ӥ��K�o��jx��\�,�I$(ҽ�B	.0��J�����A�����͎
�GL!�i�ԃA��7^��X�w�ƕO��3[��PO�p�0o�Qg�T�8��������m:��X�[�J:Jg�q�{��*�Q���8\1%�����:�aR\X!��`�v���(��!e8�baCBXBD�!�S��ZC�"�{�Q�αC]p5�N���`��٤���8���.�0uu^�aH=J�G�Dr��4N�3R���������g�W�>��̀���>�?�%�5ƥ;��2�暴���t��&��V2c+:��;*l��D�k�e-���2�]W C�;>|.��w@�ߘ5Y�K:�zQq�to�a��T���i���-ω�S�
���>a9�o���_3�|bT�M�1m���DI � �)
E�܁��u��}�*���`}�qH�i2�ys+o���U0֊`�����4n�lS�Yׇ^H�7y'Ҁ��ɼ���o��c�H~d�}C�i��=��?)���Fh���2��S�2�/��m�]�x�ރ�դ�O{:�=�|Xg�,OOO��KҞ��h��z��������s��� ��K��4�iu?��t�5N%��a�k��3��e$�vo�����ar�Ye�O��W$�2;s�or�r��-l$�s����^�N���a����OҨS1�rw%&�5v���E��y�L㥏�o含�<�w�L4`Fo'��c�����|9�Ľ �>�N���S��@KF���t�a!|F 橭�EK`ɓ�=BMe�뗶�����9h�,0�g5�܂载�X~O�<$Ѫ8����������No�E�G��4��6T�)��/M�-�t��_�h��`��k�����j��%չ�a��}κ�v��Q3�m�ܖp��"�e�T�H�A�䃯���*�o�]����B�4	nL7�8�4q���c�8��y��9i���������^������v�Ə��=�D:�I��/�y�L����w��e��L��ڦ�zqƓ^2�Y��j���D$�ϧ}v�n
��j�x-l�������&��g������%���]�7��:1t�B��������@n/e8��A�؇�Y�	><���6?m��e�L�|ǗШ�h����#���M�|�dϹ���Gh�z����Qh�$�p�sl;��(��?�ϰ��[Gԟ�E��0�c�O�K��'g����@�K��_�R0v5�Dp�y�:g��DY"�����a0ϏU҄�j�*2	k�?RF�0��[�7���7�}aS5P2>E�Fx�Z�0Y�E�7�YF�R�j7s=������x4��^U�9��M���6\ov�!99�6�"V6���W_G�� 4s+>J���i5vUf���jy�{��\�^�����JO���j��� �m~�C����K�1N)Kw�p��.Cp�����4�	d�@%]�B�H��H����aC0�����4F�`S��P���su��(W��~�0,�*q��w:�p���u�����Xe@ni�?Hܪ�O^���Pa
���]-�Cn\���sn�Xy`n +��NAU�&��V��IQxc/������^1	��le��9�UW}�Zo�G{P����4��ғ�&w���K�&�Ǚ���߷d�rR )�� ��۹=k�J�<���k�í9�w�o7P�9��e�N�=>5N.)	�^ɛ�I�5���'=����S��}���t����s1��
\	nm�$�USS+������/����o�A:� ������0�n��ן4���>�$QA���la����XU̍>⦥}�1S�A����:Ʌ����˨qH�T-��(�����+_���qc^�]��7�껔��3۲�������Y�0�
��m�9���c��AĤ��u�2���C�a�V����-+�jF-�J#�|��]%�q��~/�3uBi�@�B�دN�;������a�u_�}!��eC�X.��s�9���"�q����mT$����Ř�stTƔ�89%ߕ~�,cA��x�䃺Cb7�\}�>�ȋ��;C|WCy��X����a(�8��X��㽱 �i3� �0|9GN�=y,r�y���#%�_y"�w͜��_��
�홌H=n�ft�`�hM{�PKh�P���[�����mT{~����Y�ا�؁��g�=S��	���� :�p��	jM�f8Od��	閶�s��тd�^��s�D&�:6H>&e���
A{S#Qmb�9����.��&��I�|��Q3N�+���	7�F+D��,|��h����)��X!����UP��MX"U4
�Ɩ;�7"� �ٺ��4����oå��s�������a^��;�FK��������(��49*���K�-H��u��>���'�L�5�Di��o�#�Z��������ch�V�F}J��]�$C��?n�'c!�Qm�KB��V)Ç�z@R��{ANQD�ӄN�������KQs�������i}�$S���j}�0�{�Q���2n&���7*/i��w�SM���.oT"08H���������~�l{�(1E`�biP�֪3����i�B:�$�hf��͛0m�|�3R�ݲDc����r��� '*'�u�}X�[������NJ*�@���&N��d�R�jb<��ItRu9&"��8]�{�#P%}�K<�YM'W��N�&,D`���1�s���{aQ=�YCyV�`ֲ3�o/9"*�0F�ܯe���\� �.�����_��GhS��MM���K��1W��<�eS�����
$����'WW��
#�����\�U�wO�_4 �F��H�r�a��S�g��gsYV���\^��0R?�����U"�_�{ݮ��u*���sR�*�K8���
�
!�xR��Ѽ
&�*�/=vPƳb���&��Ui�4�*�#*
�2I����.��y*)1�cE�ж(�.��'5/E�+ֿ���7�g����0p���P@5i�ɼ|8��a�i��i�|/P��$���8
>gw�y\j��@A^�y!��)m|[70��O2��������y���q��<I%KkjG�����UF �����O�i�����ڈ��,-�
t�+*1N$r�t*Ť���%��0�~M������U�L,�l��7��X�S�CtA��?���Zda`Hu28�>���;�޳{�Z���W�9hEױ)i��SW[�����2������,��(p�����xzS���on���E��g�z��ٯ��3��%Z���