��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��r
����=o�z��5�5�����D8�Ss����q6�YL�H��Viqb[>ڒD�#�NA1���X�� �%w���h�屖��h�[��[k͘~ȏ*���Q0�s߇\��Z�����e<tl"�/�<ڼ���ϵV}�h>ک+��Z�Ӂ��2���^�C>��r����7��oŽ�cx�[khɜ�����ˬ�c�-������jr�@���t�|�JJ:z�	@ �\�Z�jP[�|�+Q��S	AA��`��T�����5��NZ�{T����E�b���<9~��E��Z���9�X�+X����]���$Y�q�#|�߾�x�tq\�[��x��}j��z�8=+d�%x3[x��-LPG�e�u�D'����1�%�f�s����C=7�e���L�xE8�L1��YR���T��73A��e����8G����2�ِU~�J���>37��r+7'��Q�M�4� ��B���/��AB���;��O��r����̠dJ��֡I

E'g�xA�������"	��ǳ���)�2�{�~�m����KPA' �]��	�1�K�:G�`7 ���u�����(��'wؾ�,���+���ocI��R��3=y��=Y$�(���ݽ0å4��>,��f �y�̀w�K[	 �]�yt��q77��b����o��`�qTm��@�Hk�1�Z���6��Fd�����ܣOq�ļ]XaH�0�
�E�I@��bE"��eJs��g`��<5{��i���'#�n|�Y쭧�{˘�wZ��_�W��$�wn,D�{�D	�ڮ�7��~"T�XfH{�E�X��Et��f�A�翿�V��D�Q��8?��[�2S��W���\�����+��[��2�d��FHiNp���90�؄U+��P��+�
Z��,�5؜m�@U.Y`��SAm�V��ۥ~#9o�,�N7�n|�.@�B5�x���b���T�k�e�b�6a�z�{��NOy]5տ�M\+�P�o�0���A=J�4��B�
4gߟ�Mi`�������T�x�`)����3~����ҩx��7�c`*X�d�?���Bx&���uH�̓��|��wRD�[��!� ^����`�b�߭�5p�dV�Ef�)�m��rf1�xX,���$lN���b]��sl��9�5n�� ����^��?W�dO�K|�fS4]�B���$7X-�\��֐^\F�5�ܶQ����i�jҝ�vv�C,��r�%��h����T�Yl�zՐ�F��ev��f�4g�����P�n�C���C.��,�ф{u)D���_��ű��}�so�{�*L�ý�^-���/�ꪄj-!@K��v���=Н6i�x�k��*}��օ��!�����M��W�����Љ��H�W8��TX�dy�Wo��w�K/\Ԡ�(lf�J��f!�yB���_k��~���N&+����{f"{��r���2��n�kx9�g�O�q�y��K��ʇ�q�d���Ƈ>���Ũ�o�9.�E�e������ox�FK������ �f�?�)ǜ�f��^����FM#�x2y�?˃*��,q3f�J@H�@X��������\��,(��W��R�����E�aX�T�{���|^͏�F���qG��g<�.��3�����%`�(���I�73�,�O$ՋaB��f���{ݾ3�w,����� ����/ ���cv{R3�)vro�u�ݠoz�^	�p�����\h�L���U|w�?�!�k|��$.�/�����c�����By��4z4ui��hn&��wK�+`�DQ �GJ�~ &!��2����֫&��`��F��|��Rz���fa���־C�K�|�����W�p	�	x�������,�P%k} a���M�g*�Y3C\���|BߺN�E~0������+!ORѮ�Y�"D�:r%��m���L��
`�Q}�r7/�'�NSe��IZ:F*���j�_b�qM6}y����&�{,�a�G^���,��B�g��k{���bi-���� B�{�o��%T��)�(�?d�R�)�׹�?غ�j&���	M$6��+�A��ZW�8������:
i����1P~�*�}?Ղ;D��!<X1�6 '�{t��ʰ����S�1�>��y�/�v���c���.C���D.����?^p�`�]t�������r��;�L�_���r"PH�.h��)k�FO�锱#�<k,c��ml"����WK�q��WI���G��g<���
�Z6�M��<w���B&H}�F��3�-)7*��}�0;����,C���V���BK�7̓�/��
����3To����M%m�
r��~ΐ��T>Gt���j"cG���v"�4t7��q�]�Sۀ;�]�ey��Lapeڿ�z$J������VZ=02J��~~V���{l=]�!�v:(%��RK�5�O���+��ak��l�ƒ���'�h�S�.0�@QX3��_�R�d����ȶ���
E��h�d��Π^��L.r��Ã��*7}�Oz�Z �H�.��5h��}<��:��W�����}�����o$�#�3��Jٞ��.�U-%Eg�S0�<��E�#���FDqV���}�ތJ��	��H�-�][K�,����F�a��qx�����|K��q�EU�$�~�d,Vj�ٙ8���<����E��{7�鏾f<�M�
i9y�4���!���?Crf��(�a�D!$��-���[We�����@zK� �����	���/F'jv0|fe���OJk3����=N��̈́�.�q2��*b9[�k�;�HTa���辒��:�и�9�aE~�H�hv�r[A����0a����/r8�ѧ�w4�/��WA������$T� .y��)hMJjD�ų�oM����ر��%�����$�2⑚3�f?�6�{����sb�i �a�"b'L[�;J�.ؖ7�s�3������ٕ���)gHIo�ɛ��G+Q��n2��B��A�8-��=/��
 M�d�9�$�	���D�T��@Mf���'����A��vӜ���*�1̱[.k~p� �c�!� �8�&�]2�='8�a%ʚ�ѳ�^�{y�9}�b�VY�9�W�y�Hå�/�6ux�z���v�x�GF��Qz��J��XO3FI�xz���z�"����P���B��|�э�=7�O�/���)��t���.�<rpx6��^�O�5��_�IH������$|M_ ��'�J��ܡf����߃���jK���H�{1�M�j1yc�O�
g��@�n�M��v��Oi���M�(����E�|��g�>T!��g��r*�;L�flKM�����h�׼C*�AjҪ�O�(
U90T��Z���ܥEO�"MP��F�?TJ������f�QA.��ᢹ������c�� �׾ҏ�Yx��gj��� m�A���c�����)�q�!i�b�5�D!*��Vf�{�n���:�)3����C�Jf�[���ZA�,o�S�����́�K,1��{��7��4:�؞����RU���Ǜ0éb�=���FB�;n	�<P�Ǚ"^-�8��GF�d���"!���[���do7'/�ݙH�.��^��[�L��;�X
�p�	���p\q�yM�7����5����I��U����Q���҈���\W&�ʏ²s�Կ�*�uyΖ=��������j�ի�+K�nh��oЇ��N���U�o��5H|p���PG�΅}١�NO��� �L#�0%Z�-2���K��P�m�"g<<�b�R�J-���x5���Cy	��]���t��b�ex>$�߶M����3�.`;yl�K����}�~bVo)��3�wL�f�Qk��'�+rȶ�X�{a�� �n���������,��՗���x��(�"N���vR���_��H���� ��%�n�.���+��Q�|KO�o�i����j�Ȁ���>�����V���tW�q{t��N�v���x�Ύ�٢թA�t�Iu����!��59��