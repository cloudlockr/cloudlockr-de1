��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�~Zڟe�tG)�Ę�Mq�Fi�B��A��P�W�l���4c�F:A�;�U������1�y��v��si����{8��  �Q�\/k�OG\��`�KdPfT�F���"�#s<j^�,ˎ�8��������77�{�	(H�y�]��]���)� ����,z���?�[|Yn���~���A<o�F�#��9o]�jx��ko�������ߞog����Bvx�Adj\m�qwJ%Bg��vu�6!����AR{WK�c�*2�0�LLP������� �Ղ�o{�;6�
�3WԴ�ir
%�L����̮>��������m����Fs)"��X���
=z�޵:.���X��W��Y�C�V��@ %��AO<;`��Bx�8x/̲0�56\ d��A t���� �y�U�o�&�@cڬ���p.r����r���;YCC�%�[�\��	o�T�ƃ�P��yZ���[��Ѳ>ȴ�UfH�
k|�)4S�l�m^�g����`���&����b���?�
�Ԅ�ʵ1�vgy�ٰ3)9n� ��#����->�~&�pR"�NB�FNZ�0n�� ���Th�a����v����/�s�@y��IcL�>&<�Xd˱-�3�j>�Um�Y�"?��>.�x)����r���(U%���U�� ʧ���#��Q��AE����x����R
a�ͪ��C�x�^�q�Ȼ���g]l��ǂR�;�p����1����e��__.*�k�B���j�n4B3Pꪧ�p���e/���E�a㓌o�5�=Y	��T�7n/�A�������K(���Q^ע(!3&����]�<�"@j�여�U�8]A=wp~ۂN���Ў��<	������>��)&n��Jx�;�6��Շ7��R�esqR�,��RGd���+��2 ��!��a�	�@��L;��RZ]A��H���E�z�l}?����������*�����M#i��5�)���[�o(wKf�Q�ڈ��=O� �S��1�@�3>�l�L�Ɔi�U)�������������5�ki�"5}��׾Tc|:���7�Y��  O�E� �|���R�cVs�	��^����US�������5����2�t�=I����`���|��	$�r9u��:��7�^ܼ���������a^gi����)t��+�o��k-�z�=M���������-ka��)b jhid��~ ��:���Y76�\�t���[���D�?w$D������F�t�59;mE��K�2qD ��T ul)ir]xvR2�|��-o����WCp}xx��ֲ����Q|�u�d�3�7����
75Rz�����^L�9�f�<%`\�P#�����<�1���3�+��Y�$�����_�}:ta_S����CLN�J�c_���#�5��s�]�Œ^ۻ���~�{A���:N.�@g+��1��j�;��S
�}P&�Q�LQ��2I�2�Ʒ,��̮�c�H�{�a�22� �	�dS���B�C��EJ���m����������\��%�FS4��u?�$ xΓ&��9ђ(������b-G�Zap,��Z��a#��+�MT���7Q#�q�T�bw й8��X�b%�+��7�c���5�=��ԑ�Z~S�x���]�e �;�'������w���r/��T.J��1��vMt�mc��?a�l?��V��/�鑛b��g�h�z��0�t�?Vc����� A�⟞��I�jn���x[�=  �s�%>�^i^�W��/�ȹ�f�9��g5	6��u��#�2/vP;I.�G���)����%�d����W�57"�^����1#� S��b���޲w��}����N�<T�P�ޔ_8�T�A,K��f��՜9"��7Z7��o�V��z��l���Jb�0��d	a��}�!a�`�	:�'Q~]v)��iR���b;�2qiRh�$}���F�c���u���v�-�F�߰�
(خ�.��+[+_t�d3�6��j��'Ї�T����4��>��Ӓ3%���s��x�%�]�8��T��p�sNF�(�Q��#m�g��bļb��>D�b�YTPi���r�L���pJo��2	dC_ �?�հ�Wg�݀"��Ε�zx�� `ř�ip�^=�v#�W���y\nh�����9Iy(�5��nG)81��u�lk�4�u#y�@r��# �um��UB�ќ�!�C��
e#'�B��j¤2D�=s"«{`�Y�!�!Mچ��%j�W��kmHܯЩ�����4�S��ù}�Qyq^o"J{'rZ�i�%òdm�E�<�5���T���mТ���$���)	�����F	����h�d���Zd��6��':F�4bz�o�
H��!C++`O��L`R�Xۅ<�4��ް@�L�36�-��\�-d�P�-�^ ���A�o���M>b~��qFh��q����?�}ytQ���D���ѐ�`�,���Ӗ�3T6�~�U�StUO�OM#��L�\
X�<۔n�f�Dřb�d������ɪ��׼���c�ۊ,�A8)j&�65���k\�I�:2��I�HAC8��k+�?�����ߑ��5���2�N�&1�t��|���SF�j��!�5��'۰��
�v�u��5ζ\TI���52�	ԤBb�=z����R���|gv�0&V��ȥH���_B�z�Ŭ�A�;��ic��i�(t�4vE8��e�p��g���+�E�z�F���|�%�q�q�;G�E��
U�_�Y/�(���5���������@v2��dY�y�Yj�6.-Utإ�9wa��n釋y��Ƒ��}&��b3w�#���e�jx�����v�Բ �_e&�<�c���wp���`��;��w	�ciY��:�lR���TA�[��Z�LqPt�V�&� ��d�@2b�6�-i��hhnTt�'���\���iOU>��􉽈�)h�+,K��ǿ;XA��~[��"*���[�+��i���P�������M���pBNm5�Q���b�{��u� Q���c7��v�ގ��:7>�Y�N"gH)�)Їc�l+;N�X��<��L���o���r��m�9T�����QP@�O8�!C��y��k
X
������5���b.ƽ����Ub����	�?�1	���2☇�}Ɣi^�9s���#�+�j�Iؙ՟�P~ɜ�˫δ�B���?��7Yj��ȬN(�=�"VPB���E��̺��9} �9$ܲD��G+��ط�O��v�p�p�����ȂOW�:��ڢW.��bO;��O�q�nu����.����(��cբ�U�oIw"����_��ӿq��7�73D������OM�k"�T�;�����
@�?��5n�^9��kJ��MJT�0@�S;��a�z����Y�{3�#{�Y���>>�[�XkL:�7�<n�5���r*�tosoz@��b����ϟx/6�"�/�G�"J~��d�ﱹ�E3CP���֜�����ZRdJ��󓌚��˾��8<�}� T�A�u7A�6D�Q���}�<����gda�^1l*bЧ�M�G�|(3��O_��|���0<K�\�kW��9�p$�g��.8��6�.礌��N��fZq7b�0�Gw��)�� уV!\ߺW$Ȼ����7���a����0��)y7�#bg�<��ojd\�#*�ӑ�f]m�F�O�����3䆚�2��^En�'L�ӎ�s����V�f�2M�p�9|�V$�������U�^֘a�zj�K��i��F�?z�se�f�=|*)�y���P�|��r7�E��b�k�-�!CmL@�IH�cu�ʃ��2k��
5����֊��,���d��xop�c�'�Oy$��Wz�������0��x��?�_wh��H��4�1�Z_('L"�>�>l^sXW�5��3~,[S��y2�OO�k��e�Ρ��t:<��7@�-flbi��ZR0��T�,��!�* �z%g$W܆q
Z{�;W��X،�>�6�\J�V,�V4ڪ�\�+
�Z'D�^*�2���J��1� x'7����o5���5����D"���B��l��p���$dM!KI�  +��H(�9��+,k�5-�o&��0:��/>)�/��&rT��lc���"�h�,Y�L$-����� /|S:w��r2c�Ǚ�d���O'=��@�JR�T��lC�_���	5�z
<��@�9u�,�Q0cU7��*��$�|�&���ީbd{���4�s�P���Qz뚙d0�>�eWc ����Ӟ
���z��8!6�i"�p\��)~����#J#�v����3��c���=�0�7�S��^ާ��j[�P��BL*��̥MK&h�U�1Uzǅ�W�x����*�L��f2�,�xd�N˚����Oj�V�$�-p��}v����xa4$�F�-�����H���Z^�N�N�<5�2���mZ��ƂW���@ȳ�yZ.��������@VRw�i\yZ�<�w+5>V��RA�I�4 �E�z�4�V���.W�tV��3���[�"��fN=)�'|�̈́a���o�\��a
���[\��/�ȶ�g	��-��yS������;����R5����G��!}�k�K����|}��t��xb݅�a��\�j�+v����4�+�sEb�1(U7�8L�Z��k�-�3�Z��
@� �愳	���_ �`�vQ��YУ����fß�0��n wVK:G��U}q]ڮ�=�.�n����DZIń9X�1�6���b�;;�IsZ\8��