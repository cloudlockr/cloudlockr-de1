��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��݊�I�W���WJ:��<�rљH�0 �\��y-X� �՝��F�j�~���F(O����L�c������
�0Omd��Rw��9�����):�D��!�j��l_�"R@k���0of��֭�J����W�\��;/&��oaX5�F�&V��]�-�6�����=#�����f��0ǡ�r� ��8ܖ����n�����>熸�.~71F/���У�}����>�{�T�a����l������ԥ��zP�F�```�Ko���B�#0����qb��~�y~��>�^;#���ww��7�`����Ch̚Z���9=>��ԇ�.�<6��.�M��Ozi�C�9ci �;�q�4�V��ީ�~r�� �tY��Ҋ�2x��	�8��B��nr��R�b��Ty��'	�%���C��F��!�}ո�#����V��qj�*`��apo�0�S��}����+�P�3@䌇)���K(8t�B�M����������=�iј�׹ry��ǅrI!���C-܁<-��s��މ����>�s-�[��iV �W�NՒ�;0������r�c!� RW{÷���ʗC�Y��F�-s)v==K��������r��s�\T�4"%��'܎���%��#rΖ+�����˙�h�QbǺ}0w�k�%U�_��2����Anr�Mȉ���dT^H2=���
��t�ϫ�ܠ�軰�bq��G�n��H��\�]:Ŵz��ԏa�ƌٓ�T�Gw��=�I��C���C4�>M/�X�ݜ}vf�y*]y'l�g�y�};�i_Q��ne�y�R�v������(��MQ�t��O�Y�fD���/;k
y�/��x��t���5��J>9g�
�C��@\Yp��J"��?����q-����*{�0��E5�=��+�^ξB4�=ao�ot��j7�����U���G}���l�㮞�Gd��>!�S#����j#\P�
��U���Bf��#$B�^>�{�A.-��sc�Tu�捃a= n�W�`�m�c��X���R&J���u����`#,�6�������wvm��f���S~��J(p/��w�GԆ}�Ƭ2[E�"�U�[�H_�4֫�K$��J�&>0Rc�F	���������F��E��<^Kyc���KpuH���($97��;�DF>$���k��	f�9���#zط ���_"��{@�G/[��k耵�g9jv��=:��Y �8F�{�z�͏�{#RIo}�L���p�_=�1JJ�"�1@pL_�5b���A�p<�O��z����: ڧy2�u|�n��E(�o��-�:�?NE��^`�\{6<�f�3�ܙje|����Rw�V�h���%Ts�P���O�0'�D�e�ޑ�ć�9$0U%/K�K��o�F��yg�7"Zg���*|F�����ؔ#�o��	��������$麖����rl ��9jA,Hx�G��o��*���]�LuE��=��Q���Q$�Bb@@%T�����$�V�ea���M�F����ɨO��� ������b����=��A��T
/?��"ޑM�P��XHn�3+UW����fl�3+�� ���Ŧ�,_2%K�u��"�)R�IX�ktɬ�
�ؘ�u`��]����Ż����/� ^�w�6[�~WU��Ϳ�ВR"d@���x��g�����$\d�1D<5��-��_2�#�،.	�`���Zz�#�:V�������"zx��ԝ=݃�}Z(1�g�{TGj��GG��L��������^0�K�����$�¨����chy��5z�{�UNF�#���8�e���L���'�P2V<�4<��J��>���g�_(QK�O>+������0<�wR���D�3��N��(Т,��d���('*(��V��s��ȅ�"]k9�)�V������.�,���r#v����P�����4Ѫ�k'�梚��t����+�<�S�k\!	B�{���%�P`as��\	(VK=�tmos����6��
LZ�#9��z�,�����~�ְ�;U2�}Aږ8e�3}+dL���k�}D|���w<
��@6��sz�h3н��Q������ׅ�[�*V�@=V-�`}�?�]�{S�Hp��łH�EN��%s��y'�3��g�;�R� ��e��<��k1�K����f��}�?����gk�����a˸ה�6��Q�Hq��8�G�z�j�(�{��2�C�t��M���Fw,�� cYb�mY%�.lV�Y���8TZ#��<�a�9�/A$u�= �ky�p6�:��Hց|��u��➔u��U1�n�^C��v�^7MD����FaXa�g�͐��='�*�¶Su�y� �u�$�kA!-z�fs����W��~H_w#� Ïe�VHƳ��<³��ס���dc]nb���l|�#��Y�;������tU�̙H��I]�qe�&�-�b��4pi�;|�ܗ�`�]����UQ�����%�}���Ei3B�2��P���IL�� `s.�,;?C_���x���#���mN��������9z����gF��5Sm��az[A���T���|�]0�͎��P�a�K�N:��f�֤y<��>ɈөF^��o�t�*,=�j�m��#���p��c�J Q唠��}i�����b��!w^L��q�y�c��]M���e�>y���C����n�i	g���W�����*)9c���#~g"B�2lq�Wa;��!2�\���v8�3�M'Ӈ�Vh�B�d�dیe-ȱJ4)������}iSً4G��4f�*i��e�^9����n�%��W�<u��P��F�x?`�B�Wՠ��)�\�N`����G�K�� ����R�+�o$���i�����C�K����c퓽��n`���֡�$\����\�D��ʊ���O��(K[��Dw+LM�Ug����R(�e$W̙��}/��G��=�q��]����5��B�9^�VK���x
�J�`��?0�:���� P�X���Tl.Ezx����G�MJ���TG��9O