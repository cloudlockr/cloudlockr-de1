��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��r
��٣�7��X=�~��'��"��z*� 9 �|4���U'k����8�)�G�����g�du��a�m
t��K�q}H?�騤�Q�(g�*Cf�1 ����Ľ�!�x���y9dZV�D33�ϖMa�_�l��v`K\���j�GE��Jgc�<`�EK���Ȇ0+�I�4�DУ�B�ΕXH<������@a0m�
J:�ؘPAǆ�.�>�Zc���n��
\�ըn�4Ӡ��R��u=���ܭB���":]������zY��1E2��h�Y��/�rC'����z���0*PHX����l`#`*��#Z=.<�c��txZQ�	�}�WcMԼ����H�����d'�k�N>���Ϻ�Ӧ!3 �)5���Βs�	@�3�ӮY8:�8��,cW#O��� ��>m��*A]Uk�1M�0~:ŀA%x�IF�y�~8�F8�K�����)#��Ү~�vg!P%���"���$��RA���bT7�.�(�lw56Ř����yX�K�e0�o��#7��Y�n5�l�^͚��V	��
���7xf�!h�F*�|5mG�%����=����w�p��P��*T��),P��u�'k�ѧO��j">:F���u퀥ttu������Zh�[�o)�<���?���C�D�.�`�������Fm���ؒ�Ep�D\��Q��4>��n�i��h=
x���S�>��Hܰ�<�͉�{.�a�Z�>���������;1e9������t�I�E�F��$xJ��y��_�����|w��
J<��ޔ����#��� ��\��\�fS�	��/%"�������H���(v�g)ðM{�>��yk��PdY&�[TE���j�\�b�@W���}��4�����R�(�,�̶��*^�:��󮿢�w��W�OqF �wT�����hkz°�/�`:���y��H4ft���=$hA3�s�\	pnM�П*)��h��s\��T�c��J.x�J�_��o�s8��~|rCV�gܑ)/;�\��3��H��� 	9Z�(��K�b�f2�қ� �g1mn���f����NK<��5�Τ���v���f�)#�X�.�$ܦ��;\�St%=A��fH����UbF���Q}-w��,O\��L"��5�E;�t���e�!���5_�V�$
�<�`|
�2w����N:���׈sg��'���rӇ�'�5ܭ���F�q֢i�X�ؼh؋��U��\τ�)��*�_��Np0�a2��9�Q9�]�`�U�4���o��Z��{�LG���+��sc��
7�>�lʃt��ҋ5�kY,�V;������{�P��a)� �A1��V�$NА��s6$7(e�I*�=�Yio�0��j0DB�9��/��5WFpwB�Z.ʤ�1˃V!X@H|����Y`_M�9<�SˬS֟L����I��s��K.�t�^>9�v��Sw�\BW�/CX�n�ē�|0�|�!��Ǡ��?��.��f���A�p�{i��'q�'����%�@"O8^�Y�)����چ����	��r�����3���RP&=��GaLk䜠�NM�B��F��}p�$j�ʻ�-��O��n,����J$0=�|�g�?�$^&���	Y��:��I��<��<����)�_�R����Snc�l�\��-йۍ)hB*�TWNϰ �\�ގ��5	%��v�u��N!��!ihky�Gۤ�������șj��<\,��G�*�Y��1�i�:\q@l���i�����Z}�7�f�gbJ_V7}���jתW��ˍ�ѱP�<O�O?���%�+�$�9�D�A_���O�pV�R�����
�F,��1������9����>�iP���� I�����