��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�~Zڟe���!Db���
�"OD���w�`�����7t�<m�l6֜s�*@����ϑ
n5Ū�/Ղ���K����� is��v�_�/�wۈj�Ȁ���gs�ȍ��{��Tf3 �^MN-�a��ь��M9S��E�������<Z�1�Ɏv9�-�-U�����U��,�پ u�"y�ꁝ-�=�q\��V���	���<$&�ef��m��3����g���C������ȮQ��BTfĎ��s�H$Dd���)��Gs\�N
Y�,��1P]o��2>v��]�B�!8a��d�����z_U��95)Sg���c5
�.@fE6�< ��;xL�E���K���`� ���^܍4r���F�g�D����(B�����!{�Ό��pv|���c1�ѕy�_���n����ȇ�sY��`b}�:�r".�r�&U�9������8�E��O��L��ujL�T�,e1a��v�����8O�ꔉ��Q[J�X 4�C7�Ot��fN���-ޢ�@��B6�0��7��vLOL�B'���'��p�.�)k_@�}�45i��)8r�!���6��d���� 9����d��BtV�����|g�\�.z��Y�&�9-Ger���1�c�����%��/���bE�өF�7�Hp��Z����M>`y�Pڰ�a7l��w��m�n�1�i�eZwfoJ��.�(j�J��[����ߐ�b��[�!��l����?�U��\Ù�ޓ�'�pΟ��=:Rź��f,[�C�Z����F�2��"��$>3��`�bNq�D��+��'|&�A��s�	M�/S�0/�ˢ�@��_} ��K�n�q
���irG��5���*1-��}�dy�ߩ�Oǡױ��G��cl������I{�^�rU������e�YЁ���4\}����7��%�����Ik���v���H�vwg:�\U$NՂ�X��U�8��g�<g��vm���mx��lY�'w�W�"&�� �!kW�_j��+"�#��ɊI�M������ņT�����m[�g
-�R{N]N)���c�4��xٝ/��� �5�����?�8�/�>�3�j��ѣ���ߑ�6��)��N{������[L�)>����Oی�o����cX�YM���%syy��b\m'4=���?\~�*�CП5;yA[=����&��T��N=�]����&d�����G��D��+�̶�tV2��H7?��QP� ��-7'����D=�l�9�+'�x:'*D����A> s%��C� \j�(��y]�U+�|����Єf#kRl�A=o�ѭ��Ɠ}��N�J�.���}f���mH�qg0kp���w�z>%B��a��,^���/��B`<L�V]A~�Ώ�2P��{�B �-�!�f�}��})@�ǃy8������-��!Kr�G׳������ڤ�\�����vA#���<����C�#����85I@�)醐#��V{�R(���j�*�qF��ը����\�(x��eu\����\��6��ٻ�q�-у�ޣHȮ$_p!��Do��7hMd v&��w0�hm��jnh�ӱmDES�7���р�6$4��r���c.Α��(4'��ܡ����7ʚ�JF���~�G�i�%NW���Di_dwN'!P߮*~ȁ���q���L��\n��J�u�Vo?Z\�����9�>����dk���Vd$�9�o�D�o�t+��P��=����^�b�j�6�\P��0����H)�LOC�rn��B$�rY���a��ւN�<8���i�4K�QR����@�����	�	Tŷ�ԟ[x�R�I���(\��m�X��n�۵ N��q��eL���$��t�E�7�t�!��:����LY���R{�Pī �:<��
{��Zk���r�2����V7W\e������j\	��H$�(t�F/w�9E	K��^\:�2�aT���恈�����#��!=��Ɩ��3v�؁]K�T��G�d�Z�2#}�&���!�dl0�&�;�^rXY؞T˟�������o�n�F'0�7��RLX�u�����QL�ʎhk���M��$_��B쒵�b��Uz{��0-�?	�g�q����̐EZ��?x�Dǂ��G�Հ�7����t�6��/�9yQ*���.[��[���4�,�`o���_"���bcTM��9dDQ�HVxC������ͰVBF�P���e�Ȃ��yi��A:v�t��i=���^�H�g�Q}��4TR�H�fҝ����/I:<3ul'kK<����R�9e�+�����<A�G	����f|`�����+R܈l��|�r��r���͍�|rF�%��#^~2����3?D���p:#��,q�Ng�N#A�xʆ&iVk,z��+�j��"��>e�5���3��S�N.�2|���