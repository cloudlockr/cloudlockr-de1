module AES();
endmodule
