��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�~Zڟe�{S߃���s,o櫨E@�F��P����C>�A���<\U5<�MV�bໟo��f�ȟ�[W�P���M������[/��Qm���\M�e��*��J���M����2P��@�2+�Uy��3�a�M�7�����=�=���0�Y�R�X=#C��Hx���1�:�,��ʻro8˜n1zE+���	 �eU�S�Kh��kQ�[�8<n*���Έ��]�md��[�E\FN){���3�ğ��F�NJ�;h� �F��6�8�9u�k�wQ��pP���ij.$W�"ɖGi�7DOѧ�{�)M��w'&�R�D�$�\�������Q���U$�[]�`�x�D��N�G ��n!���ο�|�T|f�S%Sش�\����a��v&#l���U�k��<#��ض	.����6�wYQ����7c��Q9銥��_��S&<F���ˣ����С����O���f���Um��f��*A���������T໌|9K�Q�I� ~��/L��Z�7�AF��dJ��9�wRZݟĩ������-{$K,��÷&�5�R���줌��x\.!pp-y�?�V �c����#�z�?��g��uV˧K%t7Op�k5�[Z��}�şlq�w`�����v�"g}�C&̃=�ᇗ�{ A4!�e����e��8r�}@^� 8��g�û���#B�k��	��6����
�P��ȩ�����>Cf�JL$)ֿ����s��lM���]��Ы7z���E{��`�=�s���
���ž4�]ЃJ���p.�3��R	�Sx��[�K�\U��Y$O���4���Q �f>�����m�4�%27��,e�|劗UEvVp�Է���;�w5���ݩs E&�گ0hZ�O�D!J�7���%�ce~4��K!7�j�H��45h�^2
�q� \,���9ix��].��0���/���ҡ%�6�x<Wj���߯���O���hHG�`f(%6�zH�Le��N�������guml&���oa�$�#p�E���ƿ�x_*a?��h�J���R^�<YiQp��5�̶���������E����$�Eb��*}�8��!�1�>$ݡy�}ؠy���i(X�C������ ��fXBed����jw(6��BR���d�ɉ g�w;[F�PR�(��FG+�(��\H�D;�z;�\|b�V��e��Xy?#G+�F�NI������Y VUƿ)��?Z0�W�,��z�u�. ���,��t�7�)xS������.��-d�=��	���5r����GS*��&�%�Sƨ�g��T��7�M(v�v�,��Ћ�0��Ss���Ƙ�a��P�R=!O>�5�n�g��a��E�u���ad"G������<�Z�S�PR��^���m�b��Au\���*��Q8!�#kiw�����&��f�A�b5艟�T�>�"��?�,Dmld����������~�NO<�yB\�ܳW���+�e�G�����YoVq/V0�i������^E�gh�7C=�GB�{�*�6��:G��������i5ܗ���o�D�M6N���EN�s �X��=I���Bغ,��u��!<�Xq�:G��o+�
�1M/�ԇ�*��i�����TcM��-��C[�1�u��O19��k�:�����y����V$�2���\|dᦤ��;s2,�XYڬmf�P�,�#�&8��Q��I�N+`��M�_��{�N���M�� @i>�Iÿ��MW%�j�P�Aw �7�ՅW��u�BL����㑣����Y���w�%���DS<'.�����|tQ��N�����=��b��e��w�r�繈�tU�{ClmY3��[֊$�
��v�{�"w7�,q�nA�G]���w��ݻ�O7��	�c����=�7�	��Q<����;�)/=�����)���tq�yZ�H��kW���$���'���A7[�듉����Kbi�����L�>SR� ���[����|�F�����%��]K00��	R������'W�?R~����9?-v��;�������� `wߢ~r����  z�:����Q0�"an:�S���-�(�Ɩ�hf`�k�j�0�$Q(7�<q�����D�i��� �Q��J��8��V��b��%���[��)�؇ov�����9)<8
��'f>_���.��PW�4�����mg��.�\��k�����QZ'P��� ����ȭ$VHu'�Y�@0�v{�}l�$\1/%���	�v^~t�ʽ�X6���;���  ��}8��,�R$�B%�N��7)"����yx�pr*��yn�=���Gg0�;�x~�(�ff��?4<U��1��S)b���w�J�Rzjt������v.T�9��Jl�b�R��m�@��	c�c6>.^ �eb�&�=�v��� �/�<O�]j��n��:�jOYA 53q=�ړ�N�!�b��i���w��A���~�ߕ^It���ǁ�Ò	>��GˌD�I��* ٳ\��@Pt�iZ��������4i�M,њ,�	A��{k�z���8�P�<�z�fŘԕA�cDipO��(	���G���R\��g��I��Cx;fST�t`8P�� �x��b��^�"�����<#!\~K���N|�w�ϝB}4���P��[zVo�Iʘ<���3�����s��GT�^uP���(�ͤ�z�s����Y�9��A�9���6�ք4�~ś�Ԅ�痾�?�٭���L�
'��� >���~�OM�jJ��c�G���:�/
^!���~���[ǇW�E��
�N\��ab@��Z����'u`b�).�7�(�g�3$<���<�8Ӱ"��X��r�٣v�[��}J]F��W����ˇ$�ڠX�6�v���'�Y�g����r�Zk��%d޶B���x}��J���0j�0p�4(�4�ۨ#m�`��k�)�g>�N��R-H�����|��g� ��>؋D�HR=�)+���e������ ���G7꯼�G���~W��R�d��7)G�n����W�7,g���~���v~�s���z��R?�-{��˽�|ĵ�[�RC��m�Ŏȋ�s�U��E�?��:8��铏$��ȱ�:�Y#�I�0~hAA�P�_F�Yٔ����	�ß!C"�8�5�>=�K��(J(��%�O�o�{�D8@᢮��Ū��)r���hWɖ�-�|��;��/1��^��]8=��5o�\������tY��{�z���������J�,IM��eR�4�=8��+�T��c����Lx�'c�+ڃ\��+�,�� *���hv_;G�EY:1��;V��M�!�m���,Y����6�Z���}Y���f��bL�BLE��(2������L�ҳcұ������x\�]|N����V�h�BS�%�Ǳ���T�� �y-��vP���!'S��4��E}��qn�-);:�[�wµ���I�1X�^?������/��_m��4��nD��e�
Yk�VA���&dd$u(.�~�Ļ�d�%
��y
�����T.�����K��j�Cy�d��v������Td���!����~u�� з����$YqDxG�Er�v&�p+���z.Zjg��V
R�K���ƙ�i`L8�r�L^4IEc��!=4>�Hc���N:y���f�t��Nd���n����0�2Ė����.��UO��IY��溯��Guo8��w>9�.L�曆�/�V<<���yLǘ]ކ(��j@5��A�R���\��@T�����{���;10Q�ΠF��@ejD�e�{z�;-mϐ�<���.h]���J�Lan����H{�-�C� i�u
0���
�� G*�����Ӯ65�