��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�^V�z._��>Mb4���E�R��04o���
�ͧכ�"}F��e3��
���Ch�����wɮ�Lìm�vV�wf�9���^{u�] ,c\���M�J*�GФ}�Sݛ�!�m\J�fH΢�/}Sp�<HP���˧eC��j��1PF~��`%<\ X��p��������]�;�۵d�Asp(�����>G�h�\����;��c��و�XC�f<n}c?�kj��+�S���5l�B�����e1��L~(�92�7v�#u���~�7}�s��k�a`���]�)\'�k�z�/S.ĭ�(�����O���ʼNR7�ȴ�D�C�G<�	oBe0��tɊ ��8���q)�f��#�pH�r��$re�m��f�	����-O�Sb!ʓh�_�2u	]V1vse�^���-�����3Lup)��#IXsʪЊ[��o�]v]��y�w��l2p��r�]V?�S�B�m�CYO$;����MT������@tL<B.m�M�7Vߴ"�ǭ7z@!쭶��Բ�n' "�6���&�XnҢ=��͛&G�¾��J�(�Uג�~b	*\Yp�)�� �N������]��o�=ʕ�~]�� �
�1`��e�2��p�Ԍ���j�	�����*�Sz[MK�@8�Ƣ?"�s2��v�p����vpId4TZ_�[���M�sB��R�u�