��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�^V�z._W[7��K&��9Y�He��U�&����!�J2��-Y�y ���LA^^��j!�m�<�#�a
�K@b4�� �e�$&���`b2@(ze�Z�h��Ǯ��Юg�6�~BwK�V�o�����P}�~F�iX0�T�Osg3g.x�%��e���R5��ڔ�m̩�ל6m�����o̒hd.m�$�Fi7�h���8<r��@�ͬ����W��7H���¥�2���ɢʹ�5�?���acT�|�Vq�xeE	���W�K1�\B������k�j�H�Ɯ�w�>oa��w%`嬎�PA���hH�fJ�#>�u�堖�G��me]38H�;��P����D�)B�O�B��r 7�"g�`Gǂ'�k�J{�Zʶ[�k�S?{� �������	�_��Ϳ�������G8��mK��h#��V`ÛݾK��$z�JF��9�1i�Ň2�:'#���O/��_�R��\��Z�ގO�&NH��o.�w4u�����_1�U�{2S�������-//R6�@�)�i�M��>�ǡ7S�X�	�.	a��3�G��E!U�r�ch�/����-{��-_*��kQ�܄�n��f�e�Y��r��k���N��_ȝ�ض��V�̎Y	!�B�å���%1\1�i���l��L[�����M�ː �s)3[����/�=m�6���=Qp=W�����;�"��76#���u��%I�x�}�Bb�4�|�H�;�\E
�O��;�B@WJ!�ޓ����Es`��+qU-�W�.㴰n>XuV�|�6Jj^�uL�F�7@�W���iG���P~���p@9A��s�"�z2Dݞ=t��%%�)�ܷQRԣ'������;�r�Pl��sY,�4}%����h��4��
2a-�""�:���~w՝��[����	�m����5h�w"R�i9�"[Y�R&�ܙ�z	���V�Ta���T����p��x�u��B�Szь;�n=�R�o��ޅ(P��4�B�W�"���AG���)V6E��ғ�W`5��A�/�D�%߯jW�-�m��h:�@�p�����N�9�	5�����&�BM�t�9����(��4��\�@G
Yq��b�G�$�~�A��5�-�׵F���+�@�E�Q%�v��o7[I�I�FS'R��>.�gZ�k��X#�R�!Iɰ7�<�79���z��x.���z���{��(3�Fu�����s�u[��\Us�>+�
]+�'��7R����Ύ��;8�������_�o��`Ĝ�cc16�P/X�Ǎܯ���P5�H��ԑ�&]�^����C'��4�*1yY�y�cZi6_��P�y��.����O���q2����O��L����;��v{�EnͰ!�춘OK���j�S��b�@�)�ǹҙ����`(4�϶R�~�_hd�OϘ*.�;�����P�G�=�}�����Lc-M
�#�8��?a\K�j��x%�x���
��o��Kɭ�I�LGRC\g�����_����>��[�2�5�n�����Z�t���M$g ��]�Y�o� ��6q�*��P�"���G�(�W�k���`���)K�� (eUr8b!�XT��_�p� 
Q��{	fo�[��.	Vuy��Y���'/�qy��1f����T=�6�F����J`�=c�ҋLC�×J%7��9� �]�SY��'m�z��X8�D��>�Α�i�,�_�=�|EW�瑙�I��L1m� ��D�G��,�ayŕbr>Ejg�Hqګ�V�P>E�����:~������أ�o�}�$�Y�N���Em�ɓ�1��������
���'x�������6cs�?M�Y���UW��t�A�		����G�?��b��[]i��y�z/�E}��]J��
й��L����(�M���8fl�Y�Q����s�^]��{���j�f�Z,R�Xl(��r���@���~�;�6��M�!�TN8��,4�QmZ>[�t�6�Ar�Dm=�}#�=m���I����I��oi(6�2.�oB��6sܱ����P;ܯ}�4&
��Y@X�-��(��ZG�Ǻ?����1ζ�C�e�t�������r=�]��8���<qd8�f���|���3�={JM+��n�����a�6b����X�9T�m�}��|B_N��ܼH�(c�LPk��.ۍ郁����`m:)Z�5"��f�5lV��Y_9�e���M����4*[�R /#kqiVн���2�z��b�Mp�_�?Lc�cʤ�Y>��DZlȼ���5M?�M�b�v]^+���1a�L9�k�NN�� �u�O6�3��_�9���O��	�e��5���bk���wXY����]G�5k����5K���<R����)\Z}�c�.f�q�xc��Aܿ�V�`��� x�/�s�;+��A�	��Y/��D�����4%��m�q����Sb�ܚ��M�f��C��{,n3�N�g���^Ȍ�6?'l�0nD�-��o������#��y��DSR#�e���C*��6O��ᄄ�Z�Pz���4NE�p���_NY�gJyE�h��Z��P@�M��\q-�(�&!\�|Z¦kD�R�]���P��	�֋��p�<э��:'�T��@X��oE�@y�R����thz��K�8蹶s���Z r�ns ���5<����:��Ǥ�<$4��P��Fm��ej���O�]d�ӑg[�Rk���ؕq�����H2#�z?/M^^C��*���e�^.���odp��ZE��I�}]~V$�@�tK`�Y
�/�T(p��e�@�ۊ���Z���=���kfE�G��8�*zJ��<�ϳg��1��5��'Їuppb9���&�-)��rG�|G�X,�y��7m��`:,��!���p9��ߕ��&jq�*���='�+i���$x1H�6�=ADV�@�A�-�ۤ�aJ״�o��M-���
���	֊�HO��5�B������+%�H;U��a�;iw�<�������z���FTwZ�E�z�4�֒�c.v1�co��,��R��T�=kGϨ�H%����3Ŧ��{�'���'�ȥ����n/u��<+��v��"1��5+�n'̙��M�щ�BPx)dt�i�Ԣ;d^�g��<A��]��3�|ȣ�m�sׅ��mB;2x��O��r8c��P�J3��m�ްt��M-C
l��cK6���W���
�Yr����j����@�7�Y�<*4�
�v��f��/�Y1O�^�U6��C<�����o������b�C=гU�u#c�/|��5�np�#uT�a�Y�,]d=�vNX�d^9.Q3ݯ$��bMG�b���o��Řy>�-{�����T��;�0�Vh$���Ә� �Iӗ�9�g?1[�|蜵<���h�?3���n���e$�%�J��*��Fԝa��D~p�I��2�쒛?��X����pFd��~��8�sB2�����E�=V���}Op�nb��<��f�čP�j��I��}���-2�,��52ß���?�t���+-:����&bG[5��6��u�̈�w_m�$bs]3(k�Sb�A��b�Z�0H�j�h�2���wj�T5�2^��:�QlD�Ϫ�߯����$֐@G���*\��^0$J�D��hY��6_��.�|��j2�$�z��@iO����z9T����dF�l�wf9����Ӿ�G�)�^�f���}�^y��f�D&��$��nkT�<��<`�uc̆8�XvLH��s�B����T��-�d��>9Oɳ�m"W| ��3�m�E�����q^5V5������D����� ���<� R�Rqq)��E6M]�@�}�y�W6g���-_�̯Џ��PO3J�3��o�����f�+"�r��ڞ���å�MW��nz���;�m�ȴT�ν5��E[)���x��[�P^{�ֻ[X^�{$��k$�Z�$^�o����*3��~͜�j
�pP,g�Y�u4�1�-6�7y�`H�|Bg�Op�!�"sA���WC�,}����i�B�O5�.C�$9U,��s���/��Ϸא��} O�x��-6�e�E�@D�N؃��w��
�埋Ĕ�!*R
KY�+y�?���0���io���mw��������m��{E�X�9��U�s�ЎS���E����Vo���b�� .��'I[����sKM���|�^�Y�6Nx�RtKfz��y]�!�nG+�Pr����]�b��P���>��k7�j�񆒛�޸�qZ���$�=���-L����P���t����?�Y5
h��E7'��n š���f~5CH��{�^W7�����g��,}wͫ��X�Dj�=d����m��<uJ�4�^��U�4���
S�j���<���۔�$m�����2X=ZB�WM�b'�C��Ohi�H�H�W��������9-Gviu�R34Ԥ?	�܉HS���8~�V�Fe^���+
��"Sy)zx8�5�"�@z)K��?A�5�dk&cʣ�Ho���X<<�i2�EFd�۝D�G����B|�����|��xj V{����ԭΣ�CV���Yђ�΢=�6�`�����Hz��B$�b��.뒮��=X�B��%�2��8g��W����P���5�%�U~�n�ݧ���Q��E]�8_�͔r�A����HO��q��*ڋ���O���"�������][��H�q5�����ؚ��HY�$�������p�_5�yHN�X���C�<�-�`�?�ƙh�ƩN���H�B�Βq���c��#��g��tNc��K+}�">�F��Jټ�����^�t<T��� �6s����(���9���H�û":�����EF(' F�^g�S$�:����^���v94݋T�w���"2�?+��Q���*!Δ��o��]���K�8���2�K�	���?H��0�l��U��lt���7&DN���jO�$��aTh{R��<�� *����{D��c��W˃����%�5_~�q��L䬑D�$�W��E�udwʅki(q@��j-^'n|�&X�c�b�9�g
�m�=�lHW���ߟ��M�|���H؞=����-����:@dPH�����`	���r.��ށ�����`~ٽZ��0's�O�?�.��.Ǒ����O�,z�Z������ڢ_���,b���IP�5��d��&��G����F7Z��ȏ��w��Jk.\3a���~{�3����8��Ә�|2e �
r��*����d�l�r�AG_�cW�2;>�\�'�{��G�`B�m��Q-��إ7K��8�ڡ("�Q�w��eGN��ld΄�T1�&@��?���I�W�<[����f�~�*�)�!�[�!G�[ �HZ�v��3ÞB{-��2ǄF�l����!-�/[9�(���4i��Ǧ�]�|�~�a�aB� �e�vk>Hm�7��3�1�B(�.�0'�f5������,�@p����Τ���
=r&{z�G�'��>.2A�Ja�EG.���:��T:�����J�g"���OSV��HPP�7�R��C$���{��X�ԭ���ƦnBz�3��ksw&� Yy��&SI�e�t��j���e.Y��54��vj�p���ՠ��'����F*J��>`;aN2є����@-H�L6u]�.V��y����vE��KD)������e-���d?���A��f�}0	��OT��2�� fW`5>*+ɯ�
��^S`���Ϯ��L7�kB�Q�=�كLX��g�tB�#&;
Iy��0oYK3l#)͵N��͙?m���v�C���s��F"޼X�Ȍ��x��nGn��AO�f�R��Eb���^��{�4��m
���ipP�ĳ�r	�A�S�� ~���%Q%v�'���7��4�c����=7C$l�T]�
ޖ$����Ӆ:2<)>g��yGE9�;�Ӹ�GZ/h�S�ƚ
�LǊ�6"J���$r  p2�wT�
�H��M�<���	b�p���TX�m�rw"��KaYڇ� ���'_$7��c~��(����́�GM���zM���Vi��>�ܞ�|Q���l��-VuCV�����Jt�/�a�Y�.-H5 `���"�42���<�}�䌨���Sw�+��lc5nB���ׁ��͝+*�KV�?�N��#����AU"^�����Q�Z�u�x�U�iO�����&�|q�ڦ�;`��1e8@ L�Aul�R�)Q��'�d��Od��r1��K/�M!�ݻaY����U6���,,�-:}��% đ��geĊpB��h�@���=��N-=E���"|Et70�\�4���pː�<4��$ UA�2῕U���'\k���$�X]f�w@�W^٫��Jfآ�6�3��Krr5p�D����J���
�AV`���ջ
߮Dp�o���<�{A��O%���D�zn�N�p�OZUa{�E�9�:�d�6(��!kN�OW�q�Eێ�����""Q��U��#����	�QG�5�՟�Ҽ�#,�����$!�T��!4���`�^���چm��꩓'��f��c�G�Z�j�Ƥu��ҙv��>���?Zu[<Ҽ}uR4�>�A_�'6�uI�@�����orf�T'?i9BY�����H0 f�A�/�%�n;8qf�Q��jڃ�a���[-�����h�� Jn}Ǿ`�sV��
ؑ<]S��3�C�F�XzP3�w�����YC�i��	�/	0�M�d)�1(qM��k������>c���B���I��D��]8���]�dX|�vR��z�u9���������<��}Ɣ�B/�������q�i﫝��ȩ���%EuҀi�m�/��q�+��~���˩�*�ʊ:�A���c�M*�M�m�����C�y�_�Y^(ڨ%A&0��6B���jpp&�A'S�.@�oM���ał'���Mu�|�ɀW�Ā���EW�j�dI?��K��r�b���a������j�A�6̌<��7�4���|�����:����'a?���-�|,��]�+ي���H3��`g�Ilͻ֒ �M-R�`2T�J��xbW!�i�o)'28��@��u-*�#���]�����F��F)��Y+�ޓYʽ�I2�h��#']�y��nO$fY��ʽ����f'�}�n �Ĳ����>1�n�G�B���.�D��h�4q����!r$�;�~�d1���)�:�%����H��'w�F������y�?+��TS��W��ޛBo��-�'��d�+uΡ��P�ߕM��"$^E���hQJ��bBLQ�BӌE:�K��^x��	�j�%\���f2�����
3k���r�I��e�m��w��wE�Qp���Io��RAT%�u�J���#�u����{�x2Z��K��*�k�ш5#xE(�Q�A��>X�ڷ���"�bp:��P{~��f�aF�0&�K˛\�'x��K�n0������1sR/m�M���Le��'t��#I��q=P-�#L�2��nwB� h���j�"<_���\���0t�Kf�) �W�*/Ї���^.�מ�gj[8����fHs�͏�X{�E�P�e�-֌ۊrнU\�:y�)�	IW����}��=��Y�T�U�Ŭ��y�S�ݞI ��H����d�q��8r�A]��2.���ۛk����`�x+���.�4��O�:�X����(�<�Ro"�Sk&zNQR	�H�E�x�Ͽ>�b���"��q \#e!���âO�Ot�ׅ�������?�+��i�z�¨ӑ8%������g�HJE!��O��)aR�7�T�g��>�۾R,vs"H�b���@��<�pI�Y� ,�_�E�p��)A�>f����V����C� 
��]+y���Qt Ts����PFÏ�������"�w��Z�U�b�������Oĭ�\z�b�*�;���"62@8$��7A�*hs`�2��[�A�q'��2�@򀢑Pq�]��:�5�"!-6�w�i�5�+�|�mѩ2�/���#���M�̋����N�;'���e��l�1L�::����RU��OJ���Z���3�o*�ǋ�XQ�T��=ns����l׻N�Imz��X�yGZEy�S��%2\wV�XWv��08��O	k���D���X8ٜ�cUB۷��zo�ږfU�oOs�&b�Rh1�Aw�bv2��^z�V��o�ܮ:����6$3�ۀS5rrJ��#��]39�~��[Gn�n�������pΗ	��T�^<^��?\.��� }^��������V�w�k����H��]Y#�DuT�$��/�=M�pz���,����d�y&ea�1�E��$y��~Dzr����a�s3��[���)+�7 �t�yJ��O��!�ɐ k����Q]Ulr��`Ѓ0v��3�����&k��-��H`��FK�U�����q�ekH����t���@��� �¦^��p6���|��Ŝ�1��͍��S6G
�3G��Y8�3�6�'�–�w�kut�ɇ�U� $��� s���l��-�Q�0��Wki�=>�bڛ�X�2 �J�@H<ޮF����%:ߣ%5�6{Jbaߏ߇m|�4�xԠ� ��ZU�q,H�c����F)�DW�Q��u�&�(31��o˦�5~��M�cL�L4��Ē���r[�eP��D�����q'�WF8_B������O V������^)�ʚY�MV��-ZJY%�����"��ܒb�@ċL�)���6%�F^����$/���q+�F�0�_Ƃ�	¡��B���2�uBL,�a,�v�o��9>z�������HD$`Y2��|���E��]bY�0�=r��|��`b7�k�Y� 5�9�Ika��f�g�f53̿�d��uˉ�f�H]{_4T�ktw�@��v�JѰZ3��q��Wڿ83�-a�E�ɵ�"RKL͉�*5ɹ��ǴlA�� ��Y����o�{?lk�`r��a����,z����SE��pԔ���W������>�\]���"�OFF:�t�*��9�Czx����0�t��z��-��CgF���z2�x���)��ˡ[����wEH�Mu�7�&�v�k"N�E����;sg�8����mkJO!M�*�D�Q��4πf��f.|l}��DQSU=�Nl���`�
��F|	>�vEW��c�?J�<���~r��I��t	a��x����)�CJ��k��·H��"���	��u�HAS��%¦U��9���=�cŜ����&���>ݦق�H�hs�4�{�gJ�n�?T���P2�7R��l����k��.rF��N�y5�	y1��B![Ji`ͩ��;��Ri)
V ��MB������ҹI��d��0P:q�2�Q�"Q8�r�TEX	�����W�k�[�&ء��aH$=w+j�=�҇��+�[6c%~+���]���.܀f�8���Ȥ?lhUziKznݠ@�;Dx\vz��{��t#+z-�K���f�1��ٱ��J�
F�kVE�X��k���Q qtJw��db�k��
�������^�/Vq6��#A�Qo47��ƫ�P�}����m|d��Q =޲�@�� ?mx�4`nµ�?�� ���$�޿�Vѥ�b{s�D�D���<�F2L��aB�	e����"��f�w��	�=c�[��A3��"�o�@�	v�ޒh>u7zrm���i��9�N����c���<7�����T��+�*�3G���tyH{�b��^�-��8@i$` �;��dc�$��A k��޲��X���/�E� ��c���x��� ��Xv���}T^�X��Vpt:a2�g�6�2���쫎���3�5[3�f��L���!L9�3�Y�o��h��5��o��Jl�Q�\��c��dC�l�;�����,~�is'D)D���шUl���?�>��a�W_)��ݝ ۢ��~6	���zr/��?u<�`w+�meZ8'D���]�gqu5�������e�p�����e�ac߳�A�М� � (˺t��;��O����Uv^�S�;7��bs+T �ެ0�dF����/w�a%�U�n��P8����0�h�f�';<w�q*v鋣���2�v--����_�����QR6����9S,���}��������9�������6��K��+��`�k�h�,�i�a�쭚؀�]H,@��M��JKWe��e���,_C*��w&�i��M��8U8��9פ����C
xDl�h|(VЅ���$�_�Ggk1�%̀�s�r0'�{�+��a����Y��>�����:�(?l�8x��l+LW-�U��\�3�����4�	\�!X䰗���s�4GT}O��5x�V�PX~-�LLݗ*��v��в���V���..������$�g/4����0�烃��2�d�K];�.Ս�è9��1=K�+���5���5��y�Ugl�0�Ic�O�F��GqS'����,����Z? ���������A��kiޥY��p!F�D��P�\KZ~�.�>���۹{�����'1I;�89,̜���Ȇ��Z�fJ�Ž�� O�������´�	��'s(|���ya*��xRp���7Ի
y]��.������=[s ��_�͟���j	��	���?��Aa:h�C��ӑ7�Q�X�'O!J/��Tש�|+C�
jP}9���mW����n\�J�Ɍ��uP<M0�&�+��)(!��y|�T����Z*[$�'�53����-��Zy���%��b%p$u7uR��:�[<�&In���	�+�.�{(s��	�	�T���0u�<��N�!���y�a{$�6,��p���|x��ڀa����	aR��%>�Zs2`���[��L����t�����H����L���u��;W���n����t ^Iws���u���+a˸�~�璘��(q(q�Ž^��O��X-�r�w�`O\�8��[��l����J|/�ZM+�)�������=AS��,��C�[ԖE����Pbl3�TԜ�9x�� -�V��2��A��E���s���d�q��8b^�Ӯ�~�@G���~�$PK����8Q�DV��ķ��Q#��J��ԗ�H�ȷ%=東�[�6g��CP�$da_�]]�;���ټD>�k. x��$zZ�T�45�)����ӷo�f}%��;��q�0M#���K,e���X	����jid@kW�´2�������o6Y]���Je�μ4�}bl�ʾmք݇�W�]�W�	�M��y0RyMF>2hI!���S?�e�9�m���&�3OO;�Ba�(P��?>2�<%餕�ξ���SLa6�a��H6����0.�����[g�q-Pv6i6,uhm�X��=P�G5�ߜHM�c���_Tx�<;	�����@�2~���|rNVM�\鱐��S�E�"�O�����$o��=s��&�rI�q����28[d�)�y!���l�ͬU	�нh-�����ja�Y��cc�*�4��%V�