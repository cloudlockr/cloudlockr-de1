��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��r
���X��mE�c���P�O^K�ᣗ�wE�g0� [�J��<xc��)�k)$h�9�u����=2Cj�ӴL�#��������9�%�<�Q lְ:��XYG��$��v��9*&`�g,�5O گ[����^�nZ��Z�L$[PS�����\R4"[�C�]Cc5��c��,�a�%n��g���=���&1GLIK�mz�پ6�A-�}���~��N�h��@M�^'V^C�lY��1�&�$*�~D����a��i��Z�Ԭ�F���Z a�tu�WN�E����,ʖx5�>3GT|��k�3���kv���P�\���$[糋�l+q�F� �T=+�)�3�ɽl^ �F�G���a�l�;HVRNv���~���hz s'#ܼ#߷�k�8�N��#T������4>��B}Y{���=~$�6k����#IA��^Rgr'�GL�N�yg) ſS�:ħ�7���|�y&���ʟ
B���x�m{�DV�%7�J���Wy�ٍf낟�L�qA�n�M�ngd�tqQq�o!�w�]�yG�ݏA�LNr7��_�K�_rW}h�|(�/h��vP�C�����/B�S5��[=����?>X�=~���K���T�ց����Y�t���K<M�w�P�P;�d��|����������W���$f������q���>7J|�m�Ne$)�'c%p)Uf&lޗ&8�DV'�J��SpEkzH ��0��ל�ڏi^0qFn��VT�!�l�����PdS�&s{g�#����)m�oGn*}�:[��v_�1	V����ˍ=Y�9���'��a� 
~.UC�C/��m��<.EmYFqp��
�J��h�_� f_���;��#���^�Z���a�%tK�
������
+�7䞴QG�^��>���� 
�8Y �������F(��qybЃ͚�fM(wʳ��}O.�4��M2|�oxk���J�]��K��N�g~¾�*;��X~�$�Ù<N��5�E�t.�zW��f( u-�����W������bMգ�F=P�dd�@l�7�VX>�}��2ץ�Ǫ�=�vS~�T�;�m���,Ǜ�~E��c,H�XV@~b�z����T^��ysf��؅���[X]fb�r��|>��v0�f�3����&��2��e�>6��?m��Jd��8���|ֵDmp���_ j۶�N+�7{9�6.�v(�KгS�Z@�ѫ:�`�J��B�h�D������l�U-D�g�F�D��X�%��Pg������#.����D�<D��*HG~r��H~>E��w��a�=+2��+�Nd�,�����0��u{���s�MxS{k/�{��i��}EcOb�UV�@EM�F �r5�q'EA��1�mz�X�Q����V�c_�C����>�R���gh�4�t�J�Y��P���:����霋���7�e~B|��6�Bq�y����F��p�Avvl�q>��Vɿ#� ��	���	���>y�V�+�J0�du�{�z�й�<W��K��k�;[Xҏ���5$;��Lj)�س�=7��!/��jP�>_�i�"�zX��U)���n�׍�����|�b���y0�1H�:�x��9�,}u�3�W{oy}��!h��ě�u�����L��"��,05�5<�s���DEA�N�D�YR����1谵u��� !���"D���78q>�ٻ����n?�q�-\$��E�����Q����F��@�
��y.=��J۟xܜA���f��-_��<�ѵ�6�6�5�^�N���ԏ�jE>��~g�h�Dv�`�
Ȣo��^�\u%�8�JK���v�:�B;�U�!�&���6Ⱥ�ɲ_�SOyb��{�6Į�"�9����d�z�<e��{8����e�C�H*W,��	(1%�NczhA]����Ǿd!��6���|�vA�r��Yw�#v
F��H�?˚~qɕԭ>.��,�;��~q%R��g�hOF.�Ϥ�M��擣K���Ð�w��?�����Y�!&�3�W�@�0�>O�g����7�Q����ĒA.�M�I�>���b@�#V~����GC&7k4y	M��'6~}����P�ʅ���@�5|d����c�Qԏ6%��j��i����-9�����=������5�%���/�Hr�@��sP����A
�OZm��	 �/<0���a�o�z�N���j��������mw�1�=�C��>B��u�����<aߒ����(�@��P����vj�Ӕ<�Os[��
\����{[X\�C~�u)6�jE8q����( �l&��J�"ˊ��A��'�aV��_��k�m�{��)v��ӴNJ����l�U�(q����#� ���R\(��1��=��K�>�;���������$�U����6S;�����'������_�mw�^��D�GX;/^Y���w�k2U���S�_����3�u�R� ��r|�:�I�Ct�aw*3<�1���{�عm�ν�z�A'�v+�Ov?)��9 �|�Y��p�b
WP�vȁ��h�8#n����Ȁ���*/,�D@����I��]�pe����b�J�:�2OdK ^J�Y��/��c?��lO[��1���>�*ִ�!�$��R��v~��-嚠Q6٥m�Rr�<���1��T���PE�t�`B��X$b�Mi|Yq�n��+U�#%�I@K��t좾;]W��Z��*���F�{!t�����6�]�(uo��~5��-����ܖ��l$�ֆ\��$������o�_���u��U�ZKF�;)m���,�%��?Z8����>�׭����@߿C���1		0q�A��}����Ľ��p:鈍��ix��[J����͊(`���g*rA��$5A��O�֥WOb�)�;�e#E�wx��vsQ�2%�g3�+���\q�,��ܛq��Yӭ*�������|~�҇�!��u�=+�)��m;�I>"��ts ���q�V/�N��L�d�x��zi�f3�NKf孼��I�d<��"�&�EȪ�W=l �x�whֶ��6��5P�n�_��	�Ul��Bm����qƘMt��Cx��^�&��/����jNM�7"{��W?�D�DL%�-� `�$X]y�����:J�W���6K�Յ�,�M��fc�+���r]������k��� �6�6Î�y��8�X�ܨ$76{��?�;�4��[]g��ۼ����:cc7�.n�H M���O�:YX �1�P5��a�QG��vH<IZJ�Ȼ�p��D�Ԭ�13F~�\otSk�Թd�8p^��}�GO"�b)�f:��5@�_%�f}�Y�`�QD0�*���ጼ���0���'�L۞�]���f\�Ul̬t���s��i�a�j��>�&�"�UWl"ϰ�*_��^��v�#�^c�{���2���/�I�bȻ�\���������eXh�Q�Y���V��"[B���ɞ�P��0TR�a�R�ᗌ�U��)�G�]�` b���nUyV�P�C��|��~nf꿢�P�݃�ta�wRo��aR�x�p3m��{]�����W��