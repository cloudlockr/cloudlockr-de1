��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�W8�!��?��&�~��<V��RH�+��\�p�<qx1%�:��!^�z��o2���O��֧�*�,��$8Y��<�sz����y%�b���/��缾J��@���_��R��Y�Z�j�zρ�M��cX���48���g�}y.J��j��ua2���i��xV��k�иd��68��o�Z����n{gc�Y��|��m(�������!���p�����!ܠ��_z��r��+"ɽ�o���a\+��^��,��q��+�ԍ	���n��N3Z}h.4`#�r�{"��̰'������w��ml�4� �*<z�ӏB���T$OWr��3�7��@�ړ��%��Hϭm��8W@aX��y�/��b��I2<-�D��J����u��ow�֜�G����C��H�^iV��8���ֳ��]�q�5'e��"d�N-tj`�;5�r����Hp$?��9��� �a0���IwXD����y`���~�2ݕ���A�&�c����,����N ��H?���.#a}\�f�E�ѥ8��fpc������]��u��j�X,TlC[�B��e�G=t#��0��-�Ӌ���dH�7�����QDfc��^$4|������Ky~�Z{L)�.MO���*e�w�+
9
�K���]d]�?݄f���t���Ď�?з����=s�!�Rk������M:��Ӫ�cH��w�Un(/�Ԯ�E��;�U��Գ�9�>p���GFW�;Iuh%��]flL�qp��u��T��rs9SD�h�:')U�7�՚�'�_�����ڑ�܎�X���5J2<��� >'����o��O�4.SZc���j�rA�1s���ߺǓ�Р����l;�E\l�׫��E���1�T����K�0�%�T�g�RY+Qm
����2\�~�/�$/�*��U�#QT����Hi{}��vW�@��sI��#|����%�.�!1ݛ�kR���;��[�~�S�/WL��G7���gt~:֝�`�w�Ճ}z��U�E���M�k������q�#��o�.�YЬN�$0Ej��*���Q(�R��zԋ�:�!!n+R�A�C��B��!/��re��Y��DV���pL
�C�ՉE:�&2Rk_Q��f5	#�8oiR�1���xL�zu����{Y�<BJ�w���OBYD�����Qt�+�_��Y��O˅��� �#P�L�