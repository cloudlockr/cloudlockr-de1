��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�^V�z._W[7��KAsc�S8��_5��)hfH���a���4&�k���D߯k��J�h��WN26{�v�)��}oO�i��ɨ	h�Y򟻙tLa�UO^n��V&W���i�A2[����"]*���qG,�*$�8�p���V,���q⹿�:�1X��鼗�X�D�&i�OVM��e~��'dg6P����"���Y.׀w�!ex�hK���g_���W"���KX�<�V\�M^�����C;���ð�8�����80'����<Q��=)�Q�-�dǽ~�
,����r�]��Fg4��y/n6��Kt�#�����aW�H%��҆���[|ڧ�1�n����������ު��et�%b�{.K�5E�#d[;3@կ��&�+��  �n*��"��G'��$A�e��yu��H�9���E_ƃ����}�e4���C�x��i���J���яd[�J:��������TG����R��%�����YPU��:���B�ߥ�&:��op�פ.s{#^	Y~ĩ��Z��h *˖���y�]Z�ĺY^�X:�7���X��K��
����LG����j��'�u���T�K�؅

��i�s�G+���Y��²����+ѩ,��U/���Vވ��OԔ�E��C꡸�#`�H�3ʳs8Ϣ}�sj��<��k�OL��W_��b�ܫ���K�O���k��_��qyuˋ�Ơ���D�\扟S��l��<�P������1�vX����n
�I	vt��T��qGP�'5�N:r䎇�_��2 ��yq ed��bԩ27��Ց��|r'ARr`U�5i�le:��N������wp!�����B�P���J���`c�Gn#�_���� D�:7���E�x����,`_D`�*�������R[D�U#m�^��+���S4��}�w�,��^r�}kge�S���Jj����H��_�nO��ONq�^F�ۂ��Q6?xR�'U�V�6A6`�,��.t�Dy����x���ڈC�]����L���a�C��Ҏ�� �à���<�ݞ�E��:��^���Nβ����C98�癞r��D���+�k ���91�)�|����$��Ũ�׽��jZ�5}��F�+@�E}����)^�x���~vk��)kG�ƴ�u���[)��7%�tlrS[�����:�l|P�aB���P� *��'0B��_=�fAj^�.&�7��8v̶Aj�_�&rd�!�:��>B7�.QWkͫ�	�j�bjJ�m9��qmut�)�Y��O}v �_[�X�j�X�\�������k�"ܭ�041��A*�X|�⧙}mO�>i��i�릆�Z�~D�B�kQ&��*`-F���#�A�ԇ�5R���5s�[����8 ����F�=�ОQ�kUsXPP̰V���iUɋ�6�c�Q��-������;H�W��H��@�>)��I$�0��y:��_oh�A`���b���|rg�&L�x�zvp��j�����=��O+5�����QN3��0�Hן��� ���+2�^'�ԋE����\y����y#��oZj�)s� Iø�|9��ID�Q�<�� �ꡑ��S�2YJ�f��qjk�pCp����y�R��=\};
����YP����o�5��@��	e�������;ƏHAi��t�sЯr|�����s[��x�n[?Լ }�ti�f}�*z�{ �ʝ�֡F4�O*��ؠ��$S��e��T+��x�M�����t?�Fl4�*v���X�Տ7�`̷���A`i�T��ڿ�(���A��M�gL?4���7�+.ur��oγjry\%�i=Lb�_C[Gx�$[�l��H'��g�.�������\e�����icE�����?8�F1��,��ڴ.���:�`�ݽ������b�Y�9n�\#���!8�Х�C��C
l�T7xٵ�� K�2q/q-~n�&Qg��0v�a0n�Z2���s��)�S�k~�f(��|C�L�"� �$�{u����|y]��J ���@���b[
�����}��Nd���!�A@K�2^Hb`YΌh�cV3���%�dn��e�{"ްwM�b�{�mF�����1D�<�[�ѥ2]��eBZ�|���-��o��x��Ʉ�r���$�(4�6��a���E������B�:��T��N���7�=��O�+@�sN��T��C-ǝ{�KBƖP�]k�= ʁ�7A�����hZ�Loَv��t{"��/���������`И.p| gp���
C mol�5K(�s쎧U#����|/wM�Zǔ�����:n��7�OR� �N����h"�O�(o��)/i��\[�{d2�1xG���	rW���r�D��l'�� Ab\e�B�ɂ����� ᘪh���R'��3�t%�pb=��8g���`���H;���k�Cd�K��;��G�/��dw+`� _��~0
Ti�l�3�5�,Fb��V�s"���������g���:����Dw��rVs/�g����bএ�Vy���F<KR���5?�f�s���<��iԲ;��sƨ�����]������������)����]����H"�}��e�dp�ڪ�*�����'�?}��"V�]}]�����a��
�ZOR�R.�C�T1i�C��,��\����d�ݤ��bP��tʮ�ƚ����.���?&@Wl��&~|��?$	��������Mޜ�S��k-0�i�i���Cz��ؕ�QcJ�T�A�G`3�b쑎�UΩ�PX�s��nv�O�q<6�t�hPj:�����ZK�6h����H/�2�J8g><D+&��}3�܌�+��PZ�ua�L]��I����*�d@%�&L�9�u� (�j�C�N r]eo��%7�:��SHR���������
�!B�:�B�Q9�#���@O$8��v^�c$ӛ���E�n�s�ӄȜ�"d��@7�� �p�3/�Bzma���J"�#�������H��s>#<�Ҙ���(`c�S	��Hp�ZC�;�D�x_i82�bB��r���;�yM>� Z�WK������ETs���z�|9��T���A��sֶO�n�����e4h����MuL6w���Y~G�9�˺.�2e�?�sI���0�.�F"��A/�����}5�ag�rVPD0P ��v�]��rb�+�-�36c��8p��ۉ>pB/j�?$ڈ���#K��1oum<�	7�U���=�2�ʹ���90ٔ3��\����NO����	<��~Zm�4�mV����(.}�m+%���u喣�tԻv{֏���H���V����T(�[�;�qf^��E��3��T���m#����loF0!dJƛbK
�7�ɖe�2fķ	��$�Ѽ�uadP�#n|���;ޙ-�$��
��i��y� 4-��9�2c��Ti����AK9�y=�����lZZo5f^�� �*�를���2�;��1�1U���s*�DT��g(�\�ᨵ�9��AM��\��K=����%��xV�h_���E��l4������O�UN�\����'f�btB��=��S��r��\�ul?�M��]�MI��"XI ����}�nF�hdĊ�ap��#!�xo�8�-*`�5�>���&��t���i�Q�7P�X�_�Ո�qj�.�"�h�5��~���qT2]�$]SC�U�v��ƺD���z�z�A1��;�h��4��J�	ք��B'����ڙ>q�a�e1�(�Qf%�7U����D�r���b�hoƷΗ�̣Cq]�D�1O�o>��&�=�a��²4f��}�7�̌rB��ܐ�8��I�u�_��w�wAI=|���F�$� P!�'@a*M��=/��x+����?���4.�t|կ�#�\%l�6���	�,Akx�F�M��	Jz�F�����o14��v����U=���E~��!���K�{A���ʫ:�b�db�#_b�LD��~^{��T��
$ՠ!uo�q_M���Dr�;e6� �zx�r�5���:�" ���@�h��җ�Y0IunU�k����v?I��Cب-�J�"9/g�d�X��f�����*�[N�)-����"h����M��n+���ZMҕ#۫&Ʃ�R���ϲv��$��[2R�.�,��"@����<�E���������⚆�s�*B$.�����e�������}}�Y�4���r�gc��yA�I��k�_hĹ���`8�x�{Pӫl@�>��j�,��pz(m�Uf듔7�DaG�8UČm�7Դ4T+�ڮ�K��'��#E���l�6��-�핢|��M����:=�h���Ssx��ow�.�E,;�j׬R��s�;"��f�i���M�A������9�5r��D�=�s��Q*(#�8TT�i<�yq_�Ye�t��?��5�����gW:F���@xֺv�\-D��q~Uw�Qv�rw&U�;�����>�����:c����!��D��]F�o��׾�f#I+h�I3���d�g���*�(RM�^�&�r���M���͌�n)ƒ������3r\�2�2;j���3�6�&Yb���q1nE��4����ޚ�����d	�=�N3�O�ו��֏C�C�y=�
�����4��R8+�������4�����z��%� ��@��ǻ�-	�P/Gj��y��]���ۍ�HC?A(��n�����PewZ���᪭쪾?�(�@�ՍA.J�)lXn�ñ(�r3�����fq��q2f��-��@i��u�a� 3Z��q��$�^Pe�Bߡ�1F�ek���� Z4�����}>��Y��y�� t��fͰ.�7��'�V�kZ���Y��B�cI�T�|�"t��i1��:	sJ`=캹�gڋ�ݴ44���U�G!�C#��XR���� �4]�� %Cn[T^��$�����+j	���4ʩ]��P��� }�@1�R�M-���Z��gWl���g�7�.=�ƯK)�,W8�vP��A�4UW�mA>S>�D��A2��0� ��n�c�K������13������ѾL�(݇�dF�o��4ڨ�� vF�Z+�r� ���c�
� 6n�P}[�%@'��>��~|� 	�V�ċ�G}��w81������(��\�DC����K�b�8��%yHo��2���@�u�$����8� .��(gʯoY%���JJ��TQ��{L6�)��~Xܤl�A�&�.�R�G4���;���>o�p��^��-�����89��.��Ԑ`�?�j8����(֜v�S��>�#�ff!��@~TFS��lq��kxp�P���τO ���ٍ����=�}�C2��Ȁ7�䌍�c��t«5S��S�7^=�����qp��9B�0��:0L��u�9
o�����?��̑}p"�cv�h'��I?s�Y\��<?����X��?-0�n��#�شER�:*]�E�p^�a�A��	�����X�{R�L�J��"mI�K}��nx+�x Rykt�D���s�)h����u�3�锏QBc�0�\��� ́Kh/�]9v
+!���
\u�� �	6�B��Y�Sf3�M�TbR_�l���by0�"�hTް��0��T��Vw����������0���[�T�v-̏����m�&��a�b"�I�s�ɐ�ļ/f�i�T�Jk2<�}}���u��Q�;e_ލ+0�͞[������$}f��B���~D���<��(W�կg��]�<i)�/��f����6�w`�+�׷:
����m܏�Y��h.������s]8�v_h�"ؒ���j_E�i����/��Μd�سV�-��
����J����k6��BG�)�5R*�Y�r�Rn{OFT�h�i-(]�hX��z�|��M/�tQ;e?�_����G�CgM�gE(��6�o4h
󝷰�m��%��I�+
n�E�-Ǭ�U���K����׾׼�I��B7��̝ڭ\�7U4~����<�e�ߛ�hz��T���R�/���3ZT}o���}����w(Ҭ�����BnK��Y~��+�ӾV��<�A�ks<��^@^��Ln$�f����iF���2MM�S�k� �td�t�U�!�z���P����|<���/t˪��Y~-
bSFԗ�`�qM����E���疵��pی9�a�!���3;s���0����������s%c��u�Tw�;��0{��%��&`�p4M�����7՛}�'��U��A��Ƚ<�;o���/()���S	x��"�	n��h��b�~^[��vsn0,���I"Z%�֔xZ�8���Rp�����U��9圻#��D`���ߘ��9���5'|���2�d�&���]e�B��Q�����&nx�zj��9��3'}elAW=V8�H�@�[��H�q�a�ZDH;���+���T���>�:�i'�l��3
,+Nmᶮ�Ef�����,����ڥ���_�������ԱG������>r��YW��E@�;ڶ�G���Ff�����1j��FI��� ��6O�]�i�!@��}e�.:�-����9jy����iZQJ:I|t'���%5�"���w��%z���d�o'��X���u�?A�6�{�)X�������ڲ%�f�Qj띨C�F�E��=v�tm�%��<8����[t��
�c꿙��OV�n��BZ��	\Ƅ;����l1��G�K��|f������_~0A��K"k�<�Z?(͙/H�,7u(�f�lզ��bn��?[��`Qq����4�Et�U����ۢ+1��Yj��$~�i�	��)Qu�����8(�$�?�TW<�3%��5���?���"6�!�]�C�o@��'��;KY��E�<�q��Dゐ�$�Қ���`���t-� ���%�b����� 3�O��ؼ���� �����V�u�Y��]��FYo�@�����q8x�v'�
��ph.�����S"7��3��j*mX; �`h������[���6�sg�lH��6�3�XYeS�fK�1H\�'�A���u���F%��j��(���nN�(�4$5�kobs�Ꮡe�c��t�_�4Y������2����63����;`6�󵠌;!��WA�\�z�rs%(d�g��u���ʥpe��v�ZE����6fc�
.�|�g�Ryp����pTo�Bp�9'���fn,'Pz\��zh��F�]�d���RC�<�[)ھ/�Brv�f�����;(��}+��P���XJK+����X�۹#�fm,�K�:����!����<1�>8���[�jr�Gr"��;^τVXk�A)�آ���@��hE�a�ݟ&��8ģC!CO��7��u�ҔCę�O��[R�����ș ��G��KЖ֝tE���*��S�{T["Bh4p4��M�)3Ҩ�w��.�6��Ƿ�bzq�%������V��1�W<��&@�7�/l�J'�%{ة�_��h�1RR�����0���Y���UF��R�r�ER6ī�����y��%�!�]��"�������l �{�,z([�0��%��r<������.H�z-,�k+�^���Rև�!Y����uK�؅i���L�����g�-�hf��3��l��Z�˵�'��挖����tѓI}�Ҟ������%<'԰	�zNE��'f�nGo���c-�d~�F�����J^�<�O�k\�$Dqnǌ��#���Y�