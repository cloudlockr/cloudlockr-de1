��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�^V�z._*�����͏���<CE��W�r2�0�ϊӷ8"V4������A�;�����	>�&�E�%v�OU�o�6z�A;���B��5"����ߨ����t��G�T��D��.(�R�Ն�-���p�\}�Y=��"ƻ������K��;�u���H��sCю�C.[c�~?X�����Q��+u�غ��ՙa��o*��}N����B3�K󄵉Q���ڌ��8��˭��0s,��6 �W���RU.9oXE��[׮N�e�Y�2K��@��C�3�A����Q��T]F�!-gz�<�����N���[����k�K�	�B2?�~M��}���b��r��1w��o���j��nclD�
��ep�q�0ྲྀ����tK y+"(��%�d��l��8G����g �<`&���C>�O�{#����M�B��ۘ�,j53c��l�0�˙
g;*/��X�W+AcN* � U�m�eюh�����m�*=p�
9Y�
=����]��y_t+�$�vMn�I\�Cy��rU7B!Mk
���N:�[��R 9<�L��ı����S��'��*���$
 �5X Tn_`�̌Lդ3�~,��ς*����86�����Dv�כT�WO�fO��u�7�%�]��͸��U�"GL��5��:��[rC6� c?�)W=0���{@�����(��T؝Pp���J�>��˘t��|����GBnQc����N�ɶF�l��c"�r�|�ꍯ�O9���4�m�0�Yk�#�=�"��f���9&�ͽ��&-4�����+�������� ��l���Lv�������>pzo>}�J'���\T\��:aˎ��K���Q��������{D��̣؎.2����E0�
mʽ�My��&]�P�~����F*��sb���WƧ�_�&�����|~���5�Ɠ�/���*!��HH�L?�HI��w�~��R�ӝ[�'�n�0���󚶒0�n��'7)���a&?'�q����7�0�O�o�YYr�=�u8��Ͱ�q���SX��&\�dCƤ�B?r�A+�����uL�g�3�hr0�:S����:��^�l������F5ӳ�%���#�χ,��)��P�O"Uh��]@��pY�G��{���Y�!v8v}����� ��{�|؆FW?���*��rn�]��Ѹ��l-��G�/�5�l����M�
?j�Nt�X����Ǥ�5-��A\�{1\~16i,��f&Ë����3X�F�m��̌v�.�#ߑ'��H~�T�W��:�Z/<ñCM�}
�9�y>Ff�c�fW���rS-`�3�I����C�E��,"�u~:9���/��W(&m=�Vߖ���f�io�W�#Xl��pY4P��E���"�**
��ks@�8���@\W�!����V�ehW��D� '����1=F��FgԀ�iR�&���D.��m���z��}�f��;g�όO���{�"�e�;g��ؼ��Eq�n�[����[�L�YT��pVU������x8W,S9�S+Œ{�>EZ1�K�59���:��M�}���֍Λ�?���+c���j�Ưro��5����38�v�=��z���}�\�E�5�("��,6B�[��4y�Cf2�"��:�-gy ��<�@��n�S��O�F9�_S���i�5�wtBR����Ƨ�/7*�-XN�&�Û �U���U�|(�����"B���$��}#��
�D�R`�>N���^lO�\Q_nn��Y��C����Z4'$��7����(����`����u�&ǌ���S�N�v��c�7��^fG�ى�g�t}̑��M���4s���rY�o�\�EѠKj�F ��3�:98�zL�4:l��K�àz�)�1���OViFEt�B�W&oЪ;i���oi!�E�p�����V �{�9��ۢ��C�ojı��y�8b���n�O�p������u�t�V1�υ�ܘ6�p����$�\ lv�ea�E��\��f�?�&�ށ8P����b.]O�>��ΜLV\NT�!pQU��T8��5�X��D�@���2����IE������ S����:���iPY�h��2��b�ȩk�6�x݅
�~��G)��J��sH�7o��qi`�ؿu�:�ٜ4�;�s��o����V�����ν�������O����[=������IC~�
��L��O�����]����A�~J��xoR�|�X$�����{kk�� 쒊Q�J4��m;��Z���O�,�#�:b軦��O��mƀ�T,�|va�"��TA񐡛�&����I(���AGH�DJ5Rc�y�4 �erO�mw�����q�8���ad���<���=2�.5  ��GP .tZ��Vq|3��av�o�!0����u&�*�t�<ܽ��s��	���u0����6�	�[(�p�o�N����Ɏh��Xl�����#/�dX�'����ѻ�u#�����e �PiD[}��Y+��fL�kk�p��Hq�:q�Z$�y�[.k�M�z�DV�]�E�a{ ]�W���8���o�� ���+�y���@��׏M>��۵�( !ę'��K��C��U`xL=���
ו�V3|�I��J^��ю	���瑗"6A	���aǂ��S�����q�(�E�ψkX��<Z��ƀ{�:w�l}��� )�ar6�DQ��iV������g!� (z�xȩΨ�%�IN4�N��QZ1��g��B	�$����MX��L��(^�*=�\�q�y�(�8�;�y��1��V̤�֛�.3sЇG�ĜEo���*�D}��J�N�K�����9�jsb��@yG>�]_�!=o�T��9��O���MueFhH���Y�N]{��}�����^��䭠��5�`(*0;�1?P�]�#�Y�7�Y��}�F��̮t�p[R����c�W�I���y�	C������w�%�L3@OiE���i:|���x�Fl#�#I�eG���-Eơ��*gi��_�T�p�1ըb��IEJ�������U���YL�ʒ���R��1�b��&��M��D����ށ����t3��J��ahV�cH�Bpűr���0��1<�@'`�j� ��j��� �<�eG�9U��ޛ��H��W!�fKͭ8��P���A�&|��9�_F�h�,XGS[p��R=�J<|�ؙ%���2��e�U�(��X�r_�Q+�ޛ	�9�mQ¿�O.׉����E��~��?�6��0h�!�WC_t,$�Xk�H����$����ׂ�w�%�Z�o��Яb��iϾ�c�O���"���W��<~��"[�,qeis���zs5Җ:��5��5ы��{����Fg�����n�nK�#���\Rx���[�l�����b��Uv�H��1�n��B��<[�����08�gi�XK�72���f�9���߷�ӻ)�2��V�%O8Pٚ�es�{�{-����l�j����rS4���J�%��ƹN8@k�������8����~���j�)e�iw9�ѨI�>f�����`J�@���,'P�qr�WS~�N�\��c�E��^���c>E��A�F�<����!��Ȅ��Ē6;����Lr���5�����?)�[\ ]L��Ʈ�{mW�;}j�̻������Z2|v�7�gЈS�jf��艐Ο�4 �����5�L���������I�p+�#���5�0��������bi�E�K �ڌ^�^}4��`��h����$��kM`�`��������� 絭K/� 2�y��/��`��zu+Tn~�Q߷pHw)T��K�7��
g#4���Iu����K�x�WNߥ8��/KG(�K������P���7I�|eQ,�nEh�K%ܓgl�q�Ix�$��>޴mA�b��~�c�
��)����'�[Y����g���P�%���wfm�/��D��&�p�I�r*��1�a��MFf�9Q`�s7AH�	==�S�g:�� ��,�U�����'�si\��>8b�\|��#�z9��T&S��8�[���>�Z&,��T+�0�8�}7�|��>���]������Br��cē�n�g|�o�<�q[v�]�-�/䗩s��9!{�����Bᢢ�َ4�xs����h`4elaRY�J�_o8ɷp.0@�͘�i:�c��U�/d��[f$���W���L���8�2y����\��y�T/�vӰ���#���� 5�����8}��|Rb� �!��Aw�,��uIb[;�A��6~ۤ<*%�92k9K�d�%%�#��8��07�on��՟mw�[	-�!���.��~�����[$�·��/qC�|=7�p^8 ����P9���TK��*(G��Ba�[�i߶5+!��J��=�Zu\x � *~�i�}
�P 쏮�.���d3Bn�<,:�`a�� ���'F�/F\u6l �1�_2���r��T{txV;���39�QbU��{�c(�^au������Y�My8Y���nUl�k�'�[�@��i4�i������յ���x�K'�����#G]&7I�D��gҴ�Ȓ�/'�4g��/F2O��r>�����>n�v��҈�TC;�`�iW<)��h��� j������BX���Q�h���*Ŭ
4�R0��@�)�L#��jJ��$�����/�n���|���A�m� K96w;�^���@�	F<��D��>@�'|H0��@�C5Ggw�wv�ILW�(�Y6�zҒ�D���������y�1O�nϑb�B�i	��������j&D����֖L�%F�q%&س�� 5E�`f��� -�*g}gP2,�t��|l*{�SX��=��Q�~DzJ#�&�t�j5�#���ka�Sh���d1��5y��Rw,�*��i9�%z1G@�U��W?zӇ�d}��m�ȼ7��a_�d�i�͆t��`
E9�߿���j����