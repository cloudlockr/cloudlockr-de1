��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6���t�'�%��쁻��O|]�yw�֮��(�<~;�4��%<�!���wP������� 2&wj��&r�+��>�~�J��g���8:To��Ԥ $,\�җ���L��_��ܗ�kّ�<�B�0�#@�#|o�
^��	��X��j��IWP�/��$X$(����K3��hC]���\g �Ϯr���x-��%4��is�CCfܥ�b�U2�Oa���ժ� �د];��*�p��d|���a��x�ۉ��X��Em�ah9�m1+-3Ŷg�-�o�#��b�!�K���R5���6H[�u�Lj G,<�U#��WH�m��f,�D�ɳ�C�"�$�A��N�1�ω89/��g���)���My�&�5� !����`K�5)$Xv�"���v�XMА���N��N4#4$Q�%w:l��je�%�l��#EM�E�Ț0C�}xH�Q�!EŶF݂I$t�+o�G��]}8өj.�!e'��s��J~<��r/�,L�c��{gd��.׆õ�5�Z��J����A��z��r5���d���+Ӻ�2=�O��^�G-4;6N>��SDl� ������\)Ƅ��@Kmy��=����m5�C�W�0d��(e!A9d�2$N��B�Xr�`Blp�}�ze�����*k��`&��C�"�p�N�pv���t���L�)AB���_P*�A8�+12BEg����j��;'�U�~
g�#ǯ/���'�@vZ~��v�@��gd���;�w}|+n�O�*��	M8���[s��1��ɿ��B��R ���L#�{0��=�T<y�!h0�S�AH�f�~w��/з;��J�qA�ōķ��﶑�K����wQ)_k�&�c�i�\��g��gv��M{�PP�y�y|5�Ι���oܟ�;�o0�1��b r�u��_��]L�+�����LA���4�l<�@�å<;Wq�xuv� �P;�fb�y���H�3����d�HZ�//Q��&��U1��ጽ<2K��8q�s�#�.9���w蔰a����y��+B"��R��V��K�D�]���R���5U-�/���+��0�չ=:}4�Ygc�����Z�W=A�h���nj�B+x�SA�F(GΎ����Ϊiu�ċ�{�b����NIc Ȯ.9D�ܒ��#0Y}�����n��Sº~
?ͤ,�r�l�.~~�<�����m��%����|Mr� �>0�t�ۉ|+���O��>�e@N��h�a  �k�T��`��<Fu����U�h�Gh~�'v���B��W6*ҏy`�do�]�6`��d���&"`Nm5^�_��软lmh[��U"��j!^=���kt5���.����5 R/6��r �ťW:�y>���݅�t���a-�8@|b��z�{���[�%7{79���4O\A��z+�Ƙr��ӗ�جcR��·