��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��im�T���")ԓ����Й�1P§�>�B�e�A��Ԯg����*�X��t<�~�������p��c>a`�i��4���U��[��]��b5��K>�D<eIs|l��A@�P���l�A�~u�˻��v���v����L��@�+���̡���*��&��/q�s���!w=-�|�n��U�sM��SẎ]0H� 7�u�^8�*О8�/��l��C�Y�q��;h5�r�)�����pŌT�HM䂔�_�~=��.a��l�t�<L<�טh���D�{���M���Oel]6Z�iQ��_U�A�	��ֆ�XktH�m�֧b_����D��J� z��*$:~$����sr��\�wo�L`A{J�p-�la�׷���~�O-*Y?�Ӏ�
���'ַ�ߞJe�$fx��+>����~Lg���p���ke_�{/�S)��ʚ�%o������]�!�!�ِ�i����؂<R,��������2U�ׯ�ӑJ�˹7�����R��B
)�P�~FgS�?%U˫-l*��SS7�+7=�Y��yK�P�d�[k>�}����ϟJ�6D�&��
�9a:O���B-������%ۂVs�b��76�u� ����7+���l��F	>!.��M��V8�H���@�RZ�3����r����"���Zh���A�*����z�8��E����J�u=%�;� ����������$h%2�69 �k��"��v�~ ��uP��.M>��Sω:W�oo[z�$��s�R��;h�b�~�{��n�"�������B���W��$���F��*�mv;~C����j_�tC����Z��2�M~�f��n���w������_w/&\��3d���'����9��b��{�@���桌'�!���^���Q-zm5��x6�K�$����R�����4Ҕ�E�ɷ������ذ�aIL��df��L�]w�k�wPk�Bld���� )E��Z�#�H߬�e�0�������ڛdz�*�җ�ڸ�=��y�g�}�c�#������Q��wdd��-�Ξ/ha�A/�W�'&?�E��0Sҗ������Q����!�6�"�'�-P�w}u|8�+JRS^(�q�~_�����M�y-�=e�H!�j|�y�/�o�+2�h
>�����ӷ�2�SS�}	�gP�D�W�J����D�HM|A��q�2�+'-�%���x<y�1�P4�,��;
_�AZ�Ԟ�RN���Vw�΃BGc
c�å�N�Caw�b��(�%2�H*�p���qIs��v;��̐ Զ�>���$��Ly����՞qm��d� �|�Ԩ�7jtA���Q�ws�UC�PX��3Y��`N����Zk���8i�^���Xb�����vB��w�>�{d�F����\B���6�4�-Q<����ژ�莙��M�G@Ӡ�q�>��2׎��^aBk��q�	��m��<LRP�e���V��8Qֺ�b"��ה��e��(�3'5%�둯����� �<uu�`]�%�9�2L��i#pp����+��g���L��9�oU��G���[5����x�*��v�����!�cBXM��V�]"hQJ��i�e��E^y�BM� �hb�
1���hX�+MňL8��v!�stGP����"B$ʞ����Z�ʨ��<��Ҁc�!Y���d�D� N��H��'�Eo:M������W#)U,"���U74��{��у��`��Tyoȇ�,U�k��#��#	o�7Bta��I�܁���D���[.��3�8.�h�&��D�iP�H{���(Ԭ�,�����`Vl��2w��^�Æ�$"J���5��_x?	W� Fk_B�;Ò�=<C~W8bA�8YT��U9j�~暰�&�����<����1�_	�Gh��#�s1t@����@���	m۵��\�����F��v�^N���`|t�gx����s���h�EFJж�R��]|�,H��u��Z���7�e7K����Tݸ�t!�Se�h�Ϣg#\%�&�۽U�K>
bq�~�e͗��r7�\��1y��c7Wi�Q��P�y�g9��|)�_�Àf=[ݘ���!~��A�����"ߐ־�+�/�4���Ȼ��ُ�zc`v	��\�'�K�񨐞mN'����-�cD�����0x����
kkU�㗾��'�ǃ:Z�2�Є#G=��&��1��ϻ��sG���-�6�._ٺ��bJDK��'/$�b�:C\�
B��!Pa\��3�����m�Й���؜h���)^���J	��e�S���j������[��G��pu�)�N�Lj���I{O�	�/k�����BAal8�e�����喢
^&d��0,���)c]�M:���L�_Ɓ����͋5���������&
�`mʀ�'HGV���-��#���KU7�z?�Q�C�W޿B�U���H�J� �~�R�l|WR˘g'�L��|��P�Iz ~�k�������Q�H�=�x��VZ�$Y+��.tB���#�����Ɓ�����u�S�&��D�D�͕?>W��q4�Sɔ5�=NEŘ���6{�|�n�O�[����'�������WF�+�F��"�mL�U	�lbz0kA��9&慱��3E���\D &�o�֞�4�\���xmL�9C �ƾ�0]��%τ\�0��.��T�<����F�+	���[�.��^��T{�����r���8���K����-	\/\L�=}���F�(S�N �\�Į�#���i���v"�%�R��U�g�}.a��"�#D'���g���3���@���3�i�����B�R;i6�G�Ͼ*��Z��]�x�Ԥ �]$�L�A����'4������`�4�^��y�s�n���O�T����t�-Z7��Z��Y���圁,�K�y1��%`RoKѺ2��H�W�}���k�18�~�����B�I�~m�<����W��u�4��dq���>H���zŽ
[��h��"�d�u���oJJ������x�@��*���M$
|�0��{�������^��e	Bvd!_�0	��<���F�_z�\[��ΰ�-�y���]R
u!M;�:̙Ʀo֣��8��F�d�9+��H�%)6�4��X#��B�;�
+ɹ��9�.T<��!�F>�)�^�:&N2J_�<��~�[�F�j��5��}]�(7J�y��pS<��_0n��%t���]�Of ɟ�c3fъq&�ab�g-�n3d$A2K����z4姧�J�.���Ų:�+��:G��d����'�PWp���7�s�R=��4d|m�a9A�˺�_�[��M�]�?��"����-4'P�r��>�!��Cq\�d<�ħ��Ŧ��
��?��Z;��=<�|ο