��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��im�T���vѓ}��W��-�yp%qs>`p���zr�����:̹�&bd�v��qiϣ��� ���(�<OV�@-$V���F��iG�/l�ȳ�,*Mw94a��XN��(A��x����JNAo����XM8m1Il���2�xCt�3?[F`h�P��,��@���T���P�2w��F�ǞF��y.ch�s�kK-AP�ګց�DА�ǟ�Nw�o���Rw����Tc��� N3ܮ��FH����MXX����Yf�|��~�ǯ���f�@A��V�eg�1uH�w$d�9��uQ�g���U�A�oM��L��f�q�la��8>�*V�9,7ހ�ˍ�SW.)��vH�s����U՗��cf��m���}Ȃ�F��ɞS�����5%_�[�O�"4�8��âܖ�K�̈́��5��{��D'/{��L=�o�� ����-���U�&һ^�_k"�lY�=���!��1��*/�Zk;vN}�h�����r ���61����vV�3�q�N��*>MB��BV�j�3�K��kx��˸��B8�	'�CQv��<���̃���B!���i����|���j�m)�*�	
M�2k��"��`2N��<��q�YG�4���CO�@�z�n?Ъ�<vO�EL �����g����/�>�y��)1��W9�Ay���A��wl��c󢶟ꈭ͹�H��{z�].��V]�z�RU�8:B�d����}����n��.�@I�����1q�V˦�?��K����W�F��K�*:��_��J�:�6�nF�V���B�u�������