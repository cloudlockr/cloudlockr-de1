��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��im�T���vѓ}��W�J�=_^���Z)u�;�S��˴�	Hk��H��0X9L]��$�̄4��?!������P�_��qeD��)hh}m�,|�i�ў�o�u0�����v-�ETE^8����� �T!X�4[f��@���z�=�Vl�x���U+�r�v4�����qD!}��'�.=�>q
;�٧3��Ș�W����>�����!;-��?�W��jt+٫q҄1�>/�K��U=���.�n$լʐ�o9�n�Qr^�Cj�T�aAL��"3���~��]���E�_��n�Y���=zF�xF���huL^T���󄇼�B�5��ho"(e�]�TA��iԢHP��}�IOkx�8��?kR9#��s�fH��M����~�N��6�B�ɚz�}�Ly�����Mk�g�V��FH�R�)�%E
¿�c�i�r