��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�^V�z._�６ h�M=X��m�!����a]̲6��>�Pr1G��A;�d�B�tr_q��6X%��^P,�D�'�F�(9������ĘaL�`��8Ǐ�)$!�*q7U|�p�����nGj���
b?�]z��¿�=i�塋Yw���޺��sE�Z��v���O����x��h�c?�8�i�����<��>T!Q���]�Z�Շx�Äi��o����&A;�fS<k�a2T��y���S��$DӋO�H$��l~%�z�Z|f�r$��w�{�ʘ5MCR�����}As��>��9aS6�O�А-�ً�B�J����q�_�Zk�y:�:�D�fk�@���W����̈�&��`7ʭ�2��S��:5U5(��T���֪�d�A�j�\o�oS�-h�*�Q�kH3,���XQ�E�4$��>t�w�G�9�v��I�k�:�EA�1�-��X�.��l�j��)j���	s��N@q�? �S�d*N���w&3	����ۜ��g�����t���Ȓ�8�g��T�I��������j3������<�A�(C�<�+R8x���S�X��dqG���6rx��?��=�U$�2����&�`m=z�_{�}H��&x[��2d�8�E���ӁT�,��ˬk�C�y�L�$�]\;Y��f;� �
h�O�����y^�ej%�wÞ�WI��v�'��M�ށAڥFa��E)��R�����2��!۠�( �,���(*����	�
�E��vw�'��kdt5ZY�O�%�&���PǪ�8�Z�%{S�guMD�����V/�^}�JF����>k��D��s�H�/ r�O�0@�a�[����D<����$K�_ŧ��U��9Y�ŗ����3�]��C�g�|��brLX��ĵk�z�n׬6&��<�#�p����ThFɅ��Ǟ�s�=�{�SyI���s��ģ�{�n�J0��8�q�+G>��ӕA��:��yUٞ�SN�~L�˷����K�����R��'��*`�)G�����b��6)��Q?�O��Y�Q���)���I��1d2�5���9����-e6;�r�4r ��D�da�J�� 0,���[V��P\�a\���zB?�5^ȭ}N�$�� �eh�W5�ڸ�b;.�]�_�PfRm��u��gK>$�%̞j,ax��4F���VA�@Be^�٪ʫё��-�53���^�.�)�������U$=+�^H1�QD����h۟�ȺBi��K��=�4&���a.�����!Q����.��P�B����v��3f���4o^�;$�G�L������3��V�?��q[�S��<�{A��|����#[L�w��K�V�{]��������q5�P�©��+�\�U��tJ�6�ˬK�E0�+�ك�ũ��a� �jPed�)@oԍ�n��H�Ђ���ۗ����#�����~Եq,H�;��+0B:�iI����D��)3�r2��N~c���6�q����ٴ�����k7x :���D����$�<G��F&:�-R�g�,
o��J�3�L~`�EB�D)h�~Pc�`��v�W_jj��Q���ˈ�@�ᤈ�-�:ו�hxw� �wXf���t�IL̷�npq�r�AK��4Py^<d�8���ZAx����ؠO���*���v}��n��G�l�u�P�4+��F�L)�V"��~���DMʻ�`�c�T��~�>z���=d��~���rQ�ȼH�?�zr+d���=�Aqt�9���T{G'���U|�����1	Ӌ��d+��̧���R���%7�-������a���o~�̒�ݖ�G����.3<k�gMi��v>x]D�K	;4����3�k+KԆ���A�|��	{ ���$�0BE1�rG*UGP������kӒ=��^b� ����̦n;�D��Q�/�>���L��bm�IT���%C��v'V��H{k��Q�qҷ��+/�=��1&k�ͅ������Or՝�t���i