��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�j,���Hۻ^�^���
�"�bm�p����v�O�K~���D)���u�b��Aĕ%���K����>=OC&�p�w	���3� ���ʧ����M�Zwn�5�/�����֭C0;ͥE�&ة`d���?n�f��u-F]��ߧ�s8�ú�G�.9�-������Z�_>���- |�yτ�B��4ȕ�$I�~0�7��T���(�<g�X�g%_�-��D�AM�R(FY7	�S��Gu�s��Ry�4�����~�9�|.�s�>RaQ[�����0�H[f'x����9�� �K��{I�:�o��l�y�I/�D/��]�-�)�7�^��k���,�t��k2R��'�[�1��*��,�T��7����^�*쥂�7��h��p���e�������V�0���PM>)ꅪ����'7L����S5����1�w�A��p�>$�T�Ґtb$Iet1d��W�C#Sű2���Ƣ��S�^!q���Z|��J���>�)b8\�
�:�S���{��T�R �U�a����-H�X��Y��K#y�M=e:X�$�x�RҖ�%�\Ǡ��z@�3h�6�B+��y�۹�lp
L���srg^B�i׮����	)г��q��"�L���^wW�>�5��o��Z�q��B��j�i6=