��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��r
���.������>Q���=u,#��h�9;�j�A��Jn!m�/�Z�dc�l���=�����u��$u^�;�dg#t��I�z��F�#���O s�T�gW4Ǟd��9]�pj��;��˺��՛O�	�÷�+�N��|��c.	�#8�|tt� D��yb���:E5���ڤ��9R
R� ;�@q���%c�A�D��ŉ�/�D�a��h�SP ,G������������dy�GO�M;/�ޛ��bO�Qr1�s�]���[[KJb�}4ޏ�Q��jܱf�!�o@;�|���5��Z�ҭ�"
?���@��Be�f�r���ꮐA��Х�n��<��:���4Q������i�ώ�[/ǣ/��y$�L-�}��֥�X��;�r?E��LM���S_����	����vo#"�T�:檺�:���!s�Q�q�?@V�b}��}�"Ĥ���7^/���%w�%qzR�Wx�$x�z[�˕c�#J�
��X="�XR��2�<���e�E�- ���p",>>)�KA\ˡj����	��~�N��&mEL`���|�V�.e\ƕo3r}��2s���ل f���Ĩ&�#pϾ��&�؈Z�I2q�<�g��C?�J�?ef��729�SG2�Ή�N�i4��=?���*f�"�?p2s����Icv��EP���[���jM�ǖb��F\cN\�Yb���$M��G���џ�:C�@Z����k�:�$sݽ+�𫶙|��TY���bAO���\b�R� L��"��!� �f�y�t�H5�oM��,���1�-W*B��(���~���e�nV�������^��૔ ��5���]lO���_�uh�q��4���M5x�	ﶘ���o(����� ��=��o&����#��9�^7��mU��ݖ�=b���(��0O#ۭitF�Ӱ)A�)o]:*���F)&��֦���E�<��VPz�DN~��6�"V�r� c���Lh���Z���W��o�]�J���r�� G�n-m|�I�C:	���J�g ��!y)���ج�׵`�ʎ%�_@�`���R9M�f��#'�d����!ct�F�1�~䌋(p_֚�):���1��2]�f����k��R�,�8+�/�H'u)�d�n�U#U�y�ӓ��5A<7�; 0�ݻ�>[���֙SJ�:�W����/c�6�9wϖY���Mp�m=���67X�4�(S���WH�?v;׭�L��q#� �i�f�=YZ�KJA������/ײ�P��L����͠Lfq�{C��V󻫓�3�tX�u�9��������UP4mk����?��/�~���e����O��;+��[ �w�	뱢/uA�Ny)F4���ܹLQ���*>9��4��M���IK�۹}���H��9���d�QH��A�:���CC�/��$ZM��%k$Ά_3���	W4e��q���b�	V�gbEe�3��a�.��c㝻�@��'��l
`^�)���a����f�3���n������R�k�Üw�].#@Q���#gK�K��">�[Z%@g[ѓ(��imG��r�Ҧ�[��E����#$5? �~�,M�)z��%ۘ��j�nv�o� �K;i���a�r���Z{�c�C��`�ʟ3Z���eP`7N~��EFuk�|�b�,�]W5��6���\�
.ijV�7aJ��}E�dc}'1��Q�a��c�}1�4.*��{D�y�Nb��3駨Rw��%u4�ǋ�A��G�kvvW��SÓ:��%��WH���%��z����?�Ufb��4l����P�[�a+I��=�	o����7�u�HF ms�~`iH�8��8�w�X���Cv�Zotk��w�{��N}�K2K��Wt�9�oP����_��]�&)Yn ��&��*S��^��ƃ��4�x7<Ũw�. |LO�?��J�ܒ�E�(!vϫ8$�~t��,2��ҍ'wL	3I�u��ru;�3M!�o�W�?���&`q	p��}�=�R2���Q(3�U1E@��C|	[��W�S�#R�����7��3���cD9���?y�!#B�a�{Wŀ7�䏒�tg	b�q��8��IF�'�̨���!Ş����R�����b�&��SJ�.J��5��!�����|툒�,�`W�����K/j���?��aj�X��9)Hf�]s������g�I�r� �����3҅��S�X:�� ����Z2�"k��+�DQf�%S�i���3'\�Z�\����������	����K�&@�������z�����,�}����Y�EhQǵͲ~~A�I}����$.	�5���MY���Qq�KY�B�>�0�+������p��5'C}`�Y��97�-����GHl��>���-�ʅAhaɝz����zZ�E�y;�vTpL!ze&��} ���<�ᘌs���e2��k��;"���<���sP S�ʗ���� �������zl�-l\EBV�ʿ��Jԭ��I~&�pR��̕��,��4�q"?�^_��A�5�u�_"�Ƴ��	U6h����R�vD�{c�������ļ��@����J����D�7�f�B�WU��3��r��6��'��_�'ǆ��6`����BLE��>Jd
��#���w]��P�E������qo*q��J.����p'Ow �z
���K;e]�@����l�.�����[$��>	0|Ȑؽ�!8����q��ZȂ5yC[X�(%�7U��{{~��F�	�"'�3eV�mP ]t�G�� [&f��cu��U���J>�U���L�d��8r�����C�`Cr1X�\�ZL,�� }2�x���mΎ��C�!Y� Q��+`1�bH�(Qϴ��8X:�N�� ||�
w=5��\B��#�Pg�>�%e�_ꅹQ�,%f4����hż�;�8�|[�gk��)u���u �#�R̀>�Z��y���T�pv����u�9R�? 1�P��]�.�+�]:�rc�6���J?K�TKh!s�|�.=a�_�ή�K�r�~rp���s#^u);|x(�Ű�n7��֙����[TU�a_I�	L��ط-����_��?p�? 2k;Aa�^��ggRr̦�����E�5�wܠƈ(����j=i�B�pi:P��A��UD�>2�c��vV%	ք��08�Z�*!�% ;��'��SA�QurM["�rKe�k��9�`$��vZv�KX��E��R�lΌg��Z�2��`#����$�7"�}��+Nпh�V�5U6�� L����e��O&m�����?/o��Ы�Hf��{��>k)�A$�$8��l�{���0�%i��m
=#�^-�M�� �[�hQ��=	�ʽ��@v���*���?��4Q��;���cY�S)Q�;��y�ln�s,�B!��lyڻ��?��4��q��D�t,h��7���ꋅ���v��Q�;����������F���(r�0!LWftf��l��N���g%�\�����G���#�+�t������Jm�������<��*r�@�����ˋT��쭂'�BqZ5�-i,wCP"@.g��3R�Z0�J!ߏ�Y���ی��8w�l���X[�dL��������-+���_��6,в6��<��z�N̀�eLc��� f���=\�-p^ա��(i��j�PD�hX&�CCʜ�;��rڡU!�'�_O��yH����]���(�;���h��8`ӧ��S�R�)Bd�p\�y���t����M��x��|���4����'W���)f�L�~i����$ԝ]Z@�4$�
��=$��q�B�����i�U�����2�����Rk��}�
 ٶ����ͮ�pJ�2����#���*Ŷ4s�}��*��h���Ur\q���<��>��2'��S}��`^�U�K7T]j�UH֭<_�5�8��E�� T,��m<ֶ�i����Y(+[�fE�����*3ࡋ��蝉���+q���XWW��s��	(�3�K�D!q/,qE��@�&��nH�VRy��'�4�h��m�!F;b<�r?/���h>F|0�z�I96�r��b|�!����/}�/tfn3K�g|V���W�īA714z%	kp��F������/0 u�~�fZ��h]'h�h{U�y���J]lr�]V0�!,��A���v�j*�s�0Z�.O��P��uk:Eƽ��|�T� ������鱙��ނ��ܴ��̬����v�e������e�o�A`����$l���i����<���Ɠ���>��p���N}Xl�f��"ac�9%�8����2��"Kt��\Y���)���3r��j>�"[-x���	7t%�Z����0]CC��"�����YB��v�M�Ϣ���r��C}�������-x+Y�	�kKD�`���Y�{���3O��K�n!��w�rԞ�] !dR�v���dԷ��2mU,���}ιY�s7��V;-y}���.�F@�����X�ep���4\}��K���l��}C�*~_w����ԏ�O`{N�@h¥�N�x�'�T$sy&�{��P�%5����*�GX��AE�b�Zk��j� ��`���u2�~!5g0�b�(�m��T	�z��2-:���a�O�GO&�^�ɧTΌY���
A��M���9^�o��_d��aQ�`��]N���ҧ��j�5���s."<��:�邨�mb�딶-�ݨ�PJ_�#ޑt��~��i����>V��U9�(��/�+"��M*O���2N6_IJ�9L�w��+s�֯�`����t[�wa�'��}�n�%Vhys��e;�����V��%aʑ�DWr;-g��[��	x�B�H��c�������HYD� j��XeˑV"�-:���v;�K�Z���愑x�2�k������Qljk�*��gMD���燝�Ľ�<V��R�6t��(ʛ��3#Q�I*z��Fw� Do�5ڌ��x�F��N���ά��sf�n�!�I�^��d�A N�b��r��*�����Ѣ�´�Vf�q?��7A584O�&3w����Bh`�"$Ax^l@(@8�
�L�qɘ7	����h�������r��[hb���m^���ϜCX��cg�ƪ٬#�h6�e���<����:� *���yoX�f8����[zhFڿ��ů� )ʮ��h�6����v���U/0{0^X����S�ҵ��_C�վ������(!R���F�W>����D��A2q����� ���v_DN����Z��f��$)�?{Ş��?uw�ZfL�K}��MZ��B�$��c�y�[�S f��֤�+�R��ą��1�h"���)��u�^/¥-~�̬�t����ruה5��з���[���9�<��J��knj�N�N*��T�v�r&G���h��]g��9�W����M����2��J�@Es�Z��Hd^��Σ3������A0��M-Bn�?��.	�Q�fo��T%ʰ������g��x.��|kc�����w����I�%��d,��5���1�������h%z3�$�T�h�_&����b�������E���+�����HR3�8We	f]�G#Yr8#{�_�=6��*�/lp�8���[�D�0�ؖuݓ�Vh�
����X���`1�l��LLb_���P��Y6�q�뛾�L��Z���`輡��.��l�NQg¬n�E��0>��Y7R��. ���Z��Oj4.X���JYr�[���>�E@�[����T���4� �눐x��i!�	>f����T�d��P:��1D~*������n]E��!
fƐ���C�$W��@�Û�d{ω�D�*�)sE�O6�����^�N	As˳_ͮ�<���]��C/)�6U��Ĕm�YN"��uIl��/����=�&�-�O�<��,c/5ov�U�30��o�i{�]���	tx�N\��`���H��08�����|�	��A8�b�ڮY�0������渥�K�gM�~�����O�f߁����y��y� ws��,��EF�$�!�_p��Ų���pE?�7�Ǝ���K#�~F}f$r�W�4���rҬ1�0�u����|����ڽ�g@*bZ�飋��l�� R�QP.���D��h�6A�:�`�0��f��x��uZ���3��6��<�_�b��Z	��8Gо��Qk�W��H��
����᱑+P�~V�T��MCH�P�ml �c����M�����n�d,�`w����s6�ș�=���X�D�S�q����o_;�/�M���}��wS~b)�|٭�{}�"�:*�KL��`6|���_�G�:~�EWq,�\��_��[�\�6�)��I%��Zc�۷�~������i���'�h��muפ,��lξ�2��]jߙ|��������TC���Ը��,@�j)h�*q��|C)Ē��6���|��O���Q{f+$��Փ��-ՇM��B4�X��w������*\�&e���5�(J@��m\����7lV� ��e��̖�A�K-R ې^�o��.��;ΧY�?,��{��5����q��zk#��f��n�l?�e��_ФoYJ�-����S<�讋;1�L�)j��\�Ƕ�@�C�,$������1���KX����l�j��<�BSd!�K����_��[���C:|j�X8��D(5a.�Ԯ�N^M�V�֚�߹�ֳ���;8
o^;��������JK��7>�p��.2�I)7��L������X oF�n��*�.��Hy(E d#Ii��k�ԇ�ހ���d2��y_��막��4�holT?��cX�����I�����H�Sܡ+9M?���:xd?J�A��{�c���F���I���K�����|����.&�b֗��*0f�K������~���7�T@N�'".�cy�(���a��:�p�]�l��C�ٴC�d�����no�6��xi��H<��&�5��K�)�����![�T����0��z:E���pÓR5+���M��6��ܸ�x�~]v��M�I�f 4^��Y��?�g�E螣GqRs<��;)�3 ��-�a!G��`�q�2>YnY&�0>��U74�1)���9��D�=I���Q�#R��6��GDR*��
IN����6�2�t�Lj&���tE���Տ�T�{�,(��>����/�f���T��ۊAoJjۨ��T�Tl�h��%r6d-��ο��m��R�h������]H����o���Sx�����m��i�����%h)SI��^akÃ �@z�����tZ��<Ȯx`����G���������e�L�N�Gx�/�����i�-�^�}5T\�{�6b�rB���t�S�6��/��sՁp��s0!�0�oO�*U�	��ۥ�e��d=��[�.��A��>�6rtS�D�ڦ�fl[*u��w����2j�;_���珕p����w��7~���k1�5y�S���'��8`�ƣnt�xi�h^�;��h���[�	��\v��s�A�:�tڷj����wYn��@����t��)��?��4�c]�1���������,�r�~�����H��VTC�5H��Kԝ`���c�80�-��������=�Nh�'�_c0�Vĸ)m��,9��V�E�I��0ӌ�@�i����2i����3%+�^'��À?��5��I'ǱQg�ٕ2��ßT�s��8�R�����������8=�P�B<�rB��J���5�晧�"�l'��Y;m���hAf���� �����oI����WDH��ڌ]����ո
�7�iw�f���M��B��"�g�����i)�|&m���>���&����)4��X{�]��L:فzb�5�>�y��}u��1W�칪O��Է�5TA�^��E�1���bk�,�*|�Ʒ�D
�1��zZ�3��w5�ZL@s�v���xH'�?w}��������s�����Y������=]1��)��4���Q�C�Td%ՙUY"/U�'�}r�s*@���3�Y�OZ��k壞F�5��X��rl�� �Bs+�_pȣYҞe�地���=�ٮ���}M�2�mU.����yc��Az�:m���wuz�b�??��5V�3��*;N���7���ٴeM">-�?0aq��!O©�H^%�E�]��>ɵw��P
��_^v~cJ+� �+NkW#k�Q�qt�Z��&\�Z]ЍWi���u�7�W.�~'D�fF-�]I4�
�q�,.�w��R�-
{��2����5�v�2s�hB�<ig��f�컴���u��pZsN��30����GU�׀�IE�9�����j�~�(Ն��Y�1믫����M�}g���b�!���iQQw�Ӎ���k�kL\p��)�[�U�6���"^??�őD��7Ps22汤n�,��M�nbޗZ�ԏ*��*����"��ʮ>��cY��+��w{��r������F:�Y���r��H�mhX
��lI��$��;f�o�}\���o$�L5(B�����hXpeNj�)����J=����¨��'���<Aqݑ����y�B������n�k	^6�3�h��bN���qy��?_F�ٯ9!���Ӗ!�?�'�o�#�����j�T��
�����@�2h���w��S7S$�J�o�_$'ޡ������=��{����m¬[y���x�|�#�x��f�G<j�]$�A�y�W�,��?"ɀr'v��H�s�׹��"�<�5��n<��ĩ�&I������{�4)�Yu�ӹ�j*,7���+9Wj`�V�,e��#a�ڼZ�����·�{��y��/��{�d�Y���v.��ӇPZ_T�T����K�"v�|�����Į�t]�S�6�(��9٭^���������!J��X���/��?E<�Q���2\�A�2UN}󲾩�I�d !���l�k/~�,~m�����S;�{Տ��Uy��ڡ�/O��u?��6�{q��8�Q��n�e�n(s�t �Q=³�h�a��?�o���ˊzK}o���+ f����"]}����H�7gaм���H$)�՞gz>�ɍ���F��8��Q?��m�SX�G&�@��y���4����� �t �f7�ԵهA�0;���R�"D�bq��vIG?�K�N��}b�}.��sa���PTx���5�>
�c	� �*��v7�A�)3s��9�&T��ҧu<���.$<��zg�6�F��.��N	�|���Qp[=;.Q��x�����v���?�&~�yhl����0�9�yz��o�z4�v��j��''J!�K�羿ҬQv�6�<#�'�z�424J#�V�� �!��B�]B�c`���A3�O��1������>�m[���B�AsF��2&���Ҕ^�����u��:��n�A��G�[|�ۈ��b�>��k���9U��ՙL �5%�N�k�Y�8L��-�:���wq�X{&׍����0&n\��e��g/R٧�h	��5�v	H] ��Y�g��/	�1�"E�Ƌҕj���)ʽ����ͥ�\��M�9�p�4\fA�Xќ�� ��6�9j�����-m���O�����úƀ	���*��k%E�\<��L�!x@�PXѸVy+N�J?�k[�3�ͦ��%W�D�"�8��2��F��rLiZ�=&�/�s�O���G!7�L��̀7)G@RM�l�q����+P�K�Z�|r0fZ)�*BE�9y�{�F��B=�j��
[Y���嬋L�7Z�
�BU����">�5���tA�K��lK�Qڄ�˞�T
�-�׾�x-X��{�̰��p����iF�����9���\����u�����a����!�;Q���ɒ~�v�����j�ڽd�Å#�g'FH5fk}��9����O�?@R����r��������׽Z�k�&H��0���Ʈ$���M�C��?W!�c�,G	�F��ƴ�wq��L2Qw#A
E8! Y��I'�v0�K�*��t
�G}�:o>��ȻA�2`ǯ�ƴ�{֖��u�U|s3K��a�{��8�0K/��lQ!"ʘ�*�����ch!9�J�VX��:p`L>X��ȶK���BW+��8�b_/K�_R��&zZ������f�G��X�C�H�8bGïI��yx�ߙ��Ͷu-)�b������9%�@�����@v5�)�V.f-BXY�d�i��q�'~J^��5X~������-ne��7C�����D��t�k���&/wYH�b���J(�����sVl��=�W�_�w�}oh�T'�Ȇ�}���
�����e�.T<�G,xA�h�|y)lfZ'E� ��J�H�M�6�SğZ�� �s:�,��V�s�E�s(xD4M&�@T��϶�}RF%ӗt�KeJ��S�H�{xX���1����K� O�L���y^"+�W��w��K��@���7{oE�;Ӿ54�*�0�V����>��s:�a�;0�P�,*20L��/�W�a�a�F_�kP��=�N�����m�U���-ڬ�� ��,�kP�}�ga��=�TGj}�'(���B8k�l6sGɨ8�c@����P"7����1N�N֖���0�T��m��;)�N�!���p��5�p[k67��U�|u��d���0(��O(u{�0 �\��y�g� �K��;��n'�3pa~�����P��>�ℍ�L�oP%M��:u2�3�p�IY�����Yةki[ Xe�۔>V�$����|��'@���Kh3w���T��Mj0�g�W�+��T�	�Y�!!�Z�5V��(�$/��J���D�x�Hj��R�?�
n�7=�uK��9��l�*��2��Դ&&�c�V�?�%����)�r��6�0��炶� [��0���W��wX��a�@��>%�3B�*̕�z�N=�Bѐ�x`�3�ލx����c�ޅk�у������>*|�;;}��tI�ʇ�t���(�Ŝh�tN��h"oH�9�жߪ��J��V?d�m�Q�����<O�VcZ�cf�L��d_���ui�Ǽ�U8�ZϠ��gm����D����y�����zD� ��f�=��e�|�e�u2�d�G�0�� :^1���	U����7���G�,�� Q<i��<@z���4�P�V;]��y��%X�!��%\��h;���h9͈ʄ���J2���ޭmG<�o~)p��*�Z�l�wg|�G�{4|�'���� �\&�B�$�e0�w����>t�U��PiQ�Y�I�Ŧ�{(����ȏD�x�mF>7�)��t�3��՛���n� �gh�YA��n9�h?o��l���0�,�9�aL��'q��jry)�܅'�oL��?��"�������ڬ�9Qg�y�i���)B�ޝ"~T�j^m}LHŊ@�s����)���Ν~
ͩw��<����` (3����'R����aw�	K��#�����ԑ��f!B�LD�\Y_Q6o;|��ص�b�x����[GwA{��k�o�4���+��@���M�C�{m;�Ȅ���K~�r%���	�4EQ�{�o9��*x�$s�Du�<M4@�j'�#G��