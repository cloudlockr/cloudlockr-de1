��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�_պ
V�Bx���U��T�괇���~e;)�V��$�����;s��B��%no!��7���o�TP�Sf٘"<��x���x+�d�idw�[�����+��M9"M[e�������>�c����1M����ɩ&`�A��Rn�ҌSu�i_�y�����M��V�]���rM�I����c\�����p�\:����ދq�%& ��R5��$D7
��{Лxl�'��S f"��|�����[>>�n��6����{���MK$F�
�~)�*�5|]���d���MK)DB~J��
ln��1�#�%_�{�[S|-ʉN�> 2�ƿ��ʭ<���?�eǴ�U�>����سd�"�t M���48E����Y�=C� �\�͙2E݁%󞀽��]�!��'q�-m�|*8��O-R��rߏ�g)�OJ����m��S���(%�%0�:F�'2��?�M�"+�	�Ȇ�\�{��ay�v�
���[��B���\����%��>��6љ���q�53�I��O�n��=u���\j9���dpK�S�M�!l���������W�m��4$���u���x�<���:3�2��7���3::��ly����0r��a����@ْ�O���a�'�=���z��onؖ#�zC o�ɾ�����u[����_��(!:�֣���pٳ��v��t���Ǒ�C���X�'�f���N#��ƌl=Fc"#���20!Ui�y,"H�����p2h�ה�X��X�5<Z��9��a	wM�g�~��o6�]�>�"Q��`8�Q�i#�� bڜ��,S�+�H �Dw�"I����Ot�Y�y�L��8H��~���n��*�ˑ�/q"�ĕK*5�K�"�>!v�s����v;
��կBз�l�$۱�_Hu�~qUƤ���Ӿ�P��W�����B��k�F��2ѧ9��$X��oA ����s��Ą� ���WE�b;ht���"���5�YA�`C�K��I�-�aY��cHd2r+|oV�YV;�52A�VW~�F�N@U���r�/X"`������	#�}*R��G�O�ՐS%yu�d\��4��peH\��5{ i���o�{���������0zm3�]u@�� $!�1�¼�NO��^�pEu��u�^���]�sأo� h��{TU�xX}p��$ ��6�h����Z1��9�{���|�t���j��IACd�p� �̓��Z/�;�P;6�VU�Е�KW=`wi�۬)��I
Q_e�31�����)%a?�����Lrp�j���Umd����æ�|R-�C�/K�Z@�<Qp'��A
R1��^^KU,���FDl����@�l��5�Sߺζ
PG��~o���p>�,|�"+��{1O\O�yo���4�-����� 5��Լ�g>q��dѪc	j���pU~�{���
G��z�0h�Y��n�f�$dZ�U�s����Ѿ�F1�kQ�=0l+d��I=?�f睹4�ѯ����".�IZ����]ʯ��W�����HH6�B��7��[�O�����(�K/��&��r����DhL��U�*pLr�)�g�.�����B�$�H(��&���\6��İpEJ��F�z��7�Pj�7;kody�]��Bj9����IȒEꂆ�<�^C��HT�l�ʫ��=��[���$���=�\������pD��I�Bx��ɴz
�y��Y}~4bbZm��E1nVL�YG*��B�I:�R��ж�;�(TAoh&�ό�~[��=۱�B�EWK�?['�x�5NS��5V�����ZH�G?�41�E�;�`�xE�����s���,֨�?M�����y������<Y� L�	�X�Mx+.y<��
X�4�~�a�r��%@�����.rhxnn:�z;��i�]So��?��fu