��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�^V�z._�{c��
~��F	15d�Z�<��l2�<����ǭ�6�'(aa�"W`�T���Q�L �t?A�!��e�L���H0
j<92��S��y����R9�Ȝ�,ȽR��̃��8�^��L "S��p�ax���@J	Y��P��V��=;9��D���I+lu�O�}��[�hi��Q�3�����~�,vQ���FS2(ŕ��ݚwU3z�ȣR�5���x^�L��6RR�%5� (�S�W��}�c0�4뭺�N��( ����WLS�����P��3P�e�+zJ�+�;��y���b /���� �B]@��ɗ��k��3k= �^�qa�M��~$��m�ǆ�/�(N��\��c��7e"-�0����	��S�ǀ�t*�5����C�w��<�]��J��ݡ�hE،ƮB�4v��eE�v�oF��I�{6�J5-��&�K�q��{٩�L��~�2�lJ>�I�_���1�lF2���(��o4��h���>�j �T�So`�t�9.�Nd��\b�aG)5��ų!���(�S~����}���%U���AN��V�c9J��8ѤM]���A�(�����8XE����N�"���p�KH�☇8K��Ù�OU���PH�"F��h�V �������OT��#ח=N�̫:s}��#ʘ�{��q��E�Q����I���PCI(�0S,�ԋQ��?�4�Q�wm���DWz���7P�C�N����h@�=��A!�hy&Ȅg�����@{��(&��΃���b�@��B�#�:��o�.���"�����1c�Y��x�I���͸YM|׶׉+`�V���2C�E�~	���w}���>���̲8�%u.�Ukf�M���(�)n����v׽:&�?����ɯxd/!З�㰍���A��A�;n�:�NF4��F3���EVo�P����O�@���Pc��Ӏ��֧��n��6�:�z����G���l�X3�U�C�lt��3�B.�u�V[��=�q��o$p&�����	HZv�����&c�" %��C}�=Z�Ts�@/iU��Ȯ�#|���
�KW�~�cE�8�;ɜ(=~U� ����Ak�ۖ���7�	��Ʊ���c��$�V��:R&�"0c	"#�s�����%	��im��A�������A"Q%�X�]��qVx�J�s�����-�T