��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��r
���N�	t��Ff�ה�㏓�g��a2�Ά:#\�4w������zȊ��G
6��;�Y ���Ũo��(�㍼l���Ӑ�h�E";��(����\W��1m^�ŒA���yz&�<�7[�TMk�?�jEQ�?�<��1�u��b,�Pt�?R߲�����k��;�����X��V���|�t��B�:Һ��##J��F!��[�S��.N��H���:�+B�,����gy�W\63���^�-����hh��c�e�ۏ��ph��Dԏ�Clq�ɲ�T`Ch����,���'a�L1��@����K*aߒ7!J~PXB���Np/�]�L�Z�p�Ő��"Okg�Q:�<؜T�a
kP�>����K'�>�>\���@:�
5�D+F��Ե��-?ɯ��yB��1H c��3D�j�|-�Q]?�ڌ%��y�Os��n��x6����Iy�w�>0�%�t��S��tTKAY�����^JLu6�8zp
�M�!��~&�7r#h���^��m���[��nm�9gQ��/���
�[L ^Ҡڤ��*QШQ֗���{M��4���7CT\ӕ�I@�NX�dɉ�(��X�k��$�#W�.���23`�Țͣ���H2�*�P���ʹ�C(�vm� ���L������j��Y�U���*����t��O�+]�Nb��a\6�e��H���G��P��k��@��aL�|�H�nZ6�v�Ke�?�����(�N�lQ丷�49���zW$-$�eAC
�MΝ���В�t�ᙖq����
˾0�D��Mp�2�a��V��MٷOd�(r�XU������.�����S�?�'>J��fi˝4'�/�@B�a��Y�h60�1�̗4�f���byc����1b��/�1j�Ie���lu� �hߋEf��B����l���9L]y2���U��;���xd�Yu~q(rsYj��s�y6�$���e�5ASʚ���v���x�K�Y\��rX�sR�Xˀv�횈��v�у�ݾg�Es��yu9u�`��$�-�	t��C�k�$oR�ѮRP�|S-�nwFV*p���^����Ɓ!K?�l�7��5k�����`��"�F�[�8�B@X���!��7��K����ć>�(��)��\�^�)���I
���+q�7�_��۵gjRs?�>V�e�\�2��m@�V�BiѨАg�h��!�k-��d���Lj��`�P$'tO��*rPq��/�_C�RZ%#�k����B(��М�ԐS�qâ�!���^�^�{ݫ�����뿅#��B�5���ڟ�6(�W#.k4����s��� �Q�!P�18���n���*W��k���cks,�j`���hlK}����8��Ex���|F�BE/2�x�5� C�1������\�˔}3��Sd�����5p�4�
"�w8�?؁߾����w�9�|t������8�6}��f�~�9���Y;Fo��{HS3��ܝ��:vR� �#R૩�)~���@��c���<�;��u``V�Ϡ�-�'��Ed8X���B�/L��������l�.}3i��we� 1��-;=H9��Β����"�j���~K�p����畇P�������v��Dmx�|���Қ��������o[J���*����oG�P��VῬ���ϱ���F��O�'C?|Y7����׈���3m"�8�卒����Sʰ7"��lQ��7�[�� o�Ced�)�o�	t�Y��#��@ߙ�FQ賨��۞��U��S�Aj���!py�|ࢲ�1 ��T��ؼ���+�P�pW��V�DT:G�u�)8��am����pG����0��͒���v5�?#*q3���Z���T��Fۍ;�j{�+����mw�_Ъ��8��5�D����՝�M'e���Բ�:/3�l�PX�9b|9Ik]BG,+�OWsQ����w{1]��		�Z9���z��V�>B�/#F�ݾP w��O0�?�c:ߣ���=�PN�y������oo��wxayiT�^�� uP����������u��1�>_�T���a=��C_V5��Ӕ-�>3pP��tZR�ܥ��q�|�v�Rb
�ʙ����X�k�d�X�o�6�+����5������-�y^突��a��Ƽ�7���/{F�!��=�U���rr`���ß� 	h�d˄\2$)����:�&e�oST��fU��+��� =��A��@Dl�Q�Ǝ�&-���Hƣ��;���-�W$�� ~��#R��̠~P��ؓ����e��Yzn`V;�@"I���gÎ�b��GҒ�����7E��V�e�ځY���������eU��2O��� ���LS��?�TF�Q�D��$<���kF�~?A��l'�Lg�Bh{�#��Q�sp,����ps�sZe����C\���`�mqF�CXj�>:X8QʺG՞�Z���&��B��?�
:� /o�(�4I��k�����t(�u����W ��\�0��]N�(� ��͡@ω�T9	zY�e�K �3�Z%I�W(Ǫ����,�w�h��<enrh)e��/@�^�"�)/Z�zǛ��O��������Dl���'�